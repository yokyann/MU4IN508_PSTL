-- code generated from the following source code:
--   ../RibbitVm/fail.ecl
--   ../RibbitVm/vm.ecl
--
-- with the following command:
--
--    ./eclat ../RibbitVm/fail.ecl ../RibbitVm/vm.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute1707, \$234_forever7481664\, \$234_forever7481665\, \$234_forever7481666\, \$234_forever7481667\, \$234_forever7481668\, \$234_forever7481669\, \$234_forever7481670\, \$234_forever7481671\, \$234_forever7481673\, \$234_forever7481674\, \$234_forever7481675\, \$234_forever7481676\, \$310_forever7481665\, aux7331672, aux7331677, get_int703, list_tail700, loop3732, pause_getI1712, pause_getI1716, pause_getI1724, pause_getI1734, pause_getI1738, pause_getI1742, pause_getI1746, pause_getI1771, pause_getI1776, pause_getI1785, pause_getI1789, pause_getI1809, pause_getI1813, pause_getI1823, pause_getI1827, pause_getI1833, pause_getI1845, pause_getI1870, pause_getI1875, pause_getI1884, pause_getI1888, pause_getI1908, pause_getI1912, pause_getI1922, pause_getI1926, pause_getI1932, pause_getI1944, pause_getI1948, pause_getI1962, pause_getI1966, pause_getI1976, pause_getI1980, pause_getI1984, pause_getII1713, pause_getII1717, pause_getII1725, pause_getII1735, pause_getII1739, pause_getII1743, pause_getII1747, pause_getII1772, pause_getII1777, pause_getII1786, pause_getII1790, pause_getII1810, pause_getII1814, pause_getII1824, pause_getII1828, pause_getII1834, pause_getII1846, pause_getII1871, pause_getII1876, pause_getII1885, pause_getII1889, pause_getII1909, pause_getII1913, pause_getII1923, pause_getII1927, pause_getII1933, pause_getII1945, pause_getII1949, pause_getII1963, pause_getII1967, pause_getII1977, pause_getII1981, pause_getII1985, pause_setI1730, pause_setI1750, pause_setI1757, pause_setI1761, pause_setI1765, pause_setI1796, pause_setI1803, pause_setI1818, pause_setI1849, pause_setI1856, pause_setI1860, pause_setI1864, pause_setI1895, pause_setI1902, pause_setI1917, pause_setI1952, pause_setI1957, pause_setI1972, pause_setI1988, pause_setI1995, pause_setI2002, pause_setI2009, pause_setI2016, pause_setI2020, pause_setI2024, pause_setI2028, pause_setI2032, pause_setI2036, pause_setI2040, pause_setI2044, pause_setI2048, pause_setI2052, pause_setI2056, pause_setI2060, pause_setI2064, pause_setII1731, pause_setII1751, pause_setII1758, pause_setII1762, pause_setII1766, pause_setII1797, pause_setII1804, pause_setII1819, pause_setII1850, pause_setII1857, pause_setII1861, pause_setII1865, pause_setII1896, pause_setII1903, pause_setII1918, pause_setII1953, pause_setII1958, pause_setII1973, pause_setII1989, pause_setII1996, pause_setII2003, pause_setII2010, pause_setII2017, pause_setII2021, pause_setII2025, pause_setII2029, pause_setII2033, pause_setII2037, pause_setII2041, pause_setII2045, pause_setII2049, pause_setII2053, pause_setII2057, pause_setII2061, pause_setII2065, q_wait1714, q_wait1718, q_wait1726, q_wait1732, q_wait1736, q_wait1740, q_wait1744, q_wait1748, q_wait1752, q_wait1759, q_wait1763, q_wait1767, q_wait1773, q_wait1778, q_wait1787, q_wait1791, q_wait1798, q_wait1805, q_wait1811, q_wait1815, q_wait1820, q_wait1825, q_wait1829, q_wait1835, q_wait1847, q_wait1851, q_wait1858, q_wait1862, q_wait1866, q_wait1872, q_wait1877, q_wait1886, q_wait1890, q_wait1897, q_wait1904, q_wait1910, q_wait1914, q_wait1919, q_wait1924, q_wait1928, q_wait1934, q_wait1946, q_wait1950, q_wait1954, q_wait1959, q_wait1964, q_wait1968, q_wait1974, q_wait1978, q_wait1982, q_wait1986, q_wait1990, q_wait1997, q_wait2004, q_wait2011, q_wait2018, q_wait2022, q_wait2026, q_wait2030, q_wait2034, q_wait2038, q_wait2042, q_wait2046, q_wait2050, q_wait2054, q_wait2058, q_wait2062, q_wait2066);
  signal \state\: t_state;
  type array_value_32 is array (natural range <>) of value(0 to 31);
  type array_value_108 is array (natural range <>) of value(0 to 107);
  signal arr1696 : array_value_32(0 to 8999) := (others => (others => '0'));
  signal \$arr1696_value\ : value(0 to 31);
  signal \$arr1696_ptr\ : natural range 0 to 8999;
  signal \$arr1696_ptr_write\ : natural range 0 to 8999;
  signal \$arr1696_write\ : value(0 to 31);
  signal \$arr1696_write_request\ : std_logic := '0';
  signal arr1697 : array_value_108(0 to 8999) := (others => (others => '0'));
  signal \$arr1697_value\ : value(0 to 107);
  signal \$arr1697_ptr\ : natural range 0 to 8999;
  signal \$arr1697_ptr_write\ : natural range 0 to 8999;
  signal \$arr1697_write\ : value(0 to 107);
  signal \$arr1697_write_request\ : std_logic := '0';
  signal arr1698 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1698_value\ : value(0 to 31);
  signal \$arr1698_ptr\ : natural range 0 to 0;
  signal \$arr1698_ptr_write\ : natural range 0 to 0;
  signal \$arr1698_write\ : value(0 to 31);
  signal \$arr1698_write_request\ : std_logic := '0';
  signal arr1699 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1699_value\ : value(0 to 31);
  signal \$arr1699_ptr\ : natural range 0 to 0;
  signal \$arr1699_ptr_write\ : natural range 0 to 0;
  signal \$arr1699_write\ : value(0 to 31);
  signal \$arr1699_write_request\ : std_logic := '0';
  signal arr1700 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1700_value\ : value(0 to 31);
  signal \$arr1700_ptr\ : natural range 0 to 0;
  signal \$arr1700_ptr_write\ : natural range 0 to 0;
  signal \$arr1700_write\ : value(0 to 31);
  signal \$arr1700_write_request\ : std_logic := '0';
  signal arr1701 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1701_value\ : value(0 to 31);
  signal \$arr1701_ptr\ : natural range 0 to 0;
  signal \$arr1701_ptr_write\ : natural range 0 to 0;
  signal \$arr1701_write\ : value(0 to 31);
  signal \$arr1701_write_request\ : std_logic := '0';
  signal arr1702 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1702_value\ : value(0 to 31);
  signal \$arr1702_ptr\ : natural range 0 to 0;
  signal \$arr1702_ptr_write\ : natural range 0 to 0;
  signal \$arr1702_write\ : value(0 to 31);
  signal \$arr1702_write_request\ : std_logic := '0';
  signal arr1703 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr1703_value\ : value(0 to 31);
  signal \$arr1703_ptr\ : natural range 0 to 0;
  signal \$arr1703_ptr_write\ : natural range 0 to 0;
  signal \$arr1703_write\ : value(0 to 31);
  signal \$arr1703_write_request\ : std_logic := '0';
  signal arr1704 : array_value_32(0 to 5) := (others => (others => '0'));
  signal \$arr1704_value\ : value(0 to 31);
  signal \$arr1704_ptr\ : natural range 0 to 5;
  signal \$arr1704_ptr_write\ : natural range 0 to 5;
  signal \$arr1704_write\ : value(0 to 31);
  signal \$arr1704_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1696_write_request\ = '1' then
                    arr1696(\$arr1696_ptr_write\) <= \$arr1696_write\;
                  else
                   \$arr1696_value\ <= arr1696(\$arr1696_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1697_write_request\ = '1' then
                    arr1697(\$arr1697_ptr_write\) <= \$arr1697_write\;
                  else
                   \$arr1697_value\ <= arr1697(\$arr1697_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1698_write_request\ = '1' then
                    arr1698(\$arr1698_ptr_write\) <= \$arr1698_write\;
                  else
                   \$arr1698_value\ <= arr1698(\$arr1698_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1699_write_request\ = '1' then
                    arr1699(\$arr1699_ptr_write\) <= \$arr1699_write\;
                  else
                   \$arr1699_value\ <= arr1699(\$arr1699_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1700_write_request\ = '1' then
                    arr1700(\$arr1700_ptr_write\) <= \$arr1700_write\;
                  else
                   \$arr1700_value\ <= arr1700(\$arr1700_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1701_write_request\ = '1' then
                    arr1701(\$arr1701_ptr_write\) <= \$arr1701_write\;
                  else
                   \$arr1701_value\ <= arr1701(\$arr1701_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1702_write_request\ = '1' then
                    arr1702(\$arr1702_ptr_write\) <= \$arr1702_write\;
                  else
                   \$arr1702_value\ <= arr1702(\$arr1702_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1703_write_request\ = '1' then
                    arr1703(\$arr1703_ptr_write\) <= \$arr1703_write\;
                  else
                   \$arr1703_value\ <= arr1703(\$arr1703_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1704_write_request\ = '1' then
                    arr1704(\$arr1704_ptr_write\) <= \$arr1704_write\;
                  else
                   \$arr1704_value\ <= arr1704(\$arr1704_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$v1722\, \$v1938\, \$v1839\, \$v1936\, \$v105\, \$v1837\, 
               \$266\, \$v1942\, \$v1881\, \$v1710\, \$v148\, \$v1782\, 
               \$v1843\ : value(0 to 35) := (others => '0');
      variable \$v125\, \$274\, \$v113\, \$v110\, \$292\, \$v116\, 
               list_tail700_arg, \$v145\, \$283\, \$v130\, \$v186\, \$326\, 
               \$v181\, \$268\ : value(0 to 63) := (others => '0');
      variable \$v1882\, \$v1939\, \$v1840\, \$v1723\, \$v1844\, \$v1838\, 
               \$v1711\, \$v1943\, \$v1783\, \$v1937\ : value(0 to 3) := (others => '0');
      variable \$v1961\, \$v1764\, \$v1836\, \$v1960\, \$v2031\, \$v1906\, 
               rdy1706, \$v1998\, \$v2023\, \$v1780\, \$v1852\, \$v2063\, 
               \$v2027\, \$v1733\, \$v1921\, \$v1779\, \$v146\, \$v1760\, 
               \$v1863\, \$v1812\, \$303\, \$v1830\, \$v2047\, \$v1728\, 
               \$v1887\, \$v1879\, \$v1971\, \$v2012\, \$v1947\, \$v1969\, 
               \$v2005\, \$v1822\, \$v1975\, \$v1987\, \$v1745\, \$v1808\, 
               \$v1841\, \$v2039\, \$v1955\, \$v1915\, \$v1753\, \$v1898\, 
               result1705, \$v1891\, \$v1940\, \$v1727\, \$v1799\, \$v1788\, 
               \$v2055\, \$v1867\, \$v1929\, \$v1807\, \$v1774\, \$264\, 
               \$v1741\, \$v1951\, \$v1719\, \$v1911\, \$v1935\, \$v1768\, 
               \$v1983\, \$v158\, \$v1991\, \$v1792\, \$v2067\, \$v1715\, 
               \$v1878\, \$v1749\, \$v1859\, \$v1848\, \$v1925\, \$v1826\, 
               \$v1821\, \$v1970\, \$v2051\, \$v2019\, \$v2059\, \$v1979\, 
               \$v1905\, \$v1737\, \$v1775\, \$v1729\, \$v2035\, \$v106\, 
               \$v1720\, \$v1806\, \$v1816\, \$v2043\, \$v1907\, \$v1874\, 
               \$v1965\, \$v1920\, \$v1873\ : value(0 to 0) := (others => '0');
      variable aux7331677_arg, aux7331672_arg, \$v163\ : value(0 to 139) := (others => '0');
      variable \$v151\, \$v161\, \$265\, \$v170\, \$297\, \$v107\, \$v104\, 
               \$v1641\ : value(0 to 107) := (others => '0');
      variable \$v2006\, \$87_i\, \$259_x\, \$84_i\, \$v1755\, \$76_x\, 
               \$305_i\, \$287\, \$v1916\, \$v124\, \$99_x\, \$v1831\, 
               \$v199\, len, \$v1784\, \$279_i\, \$v112\, \$v2000\, \$v2008\, 
               \$v1832\, \$286\, \$270_i\, \$101_x\, \$v1769\, \$v1900\, 
               \$v111\, \$v1770\, \$v1794\, \$v1802\, \$v2001\, \$296\, 
               \$v179\, \$v1801\, \$v1992\, \$v114\, \$v1721\, \$v1842\, 
               \$325\, \$v1892\, \$81_i\, \$v1899\, \$v198\, 
               aux7331677_result, \$222_i\, \$v129\, \$71_x\, \$267\, 
               \$288_i\, \$324_c\, \$89_i\, loop3732_arg, \$v1708\, 
               get_int703_arg, \$v2013\, \$v1855\, \$v1941\, \$v1956\, 
               aux7331672_result, \$v1853\, \$v1868\, \$327\, \$v1795\, 
               \$v180\, \$v184\, \$v1756\, \$v123\, \$v1754\, \$v185\, 
               \$v1869\, \$v2014\, \$v115\, \$v1854\, \$v108\, \$v1994\, 
               \$v1709\, \$v147\, \$v1993\, \$220_i\, \$v2015\, \$v1880\, 
               \$v1893\, \$74_i\, \$v1930\, \$269\, \$v1817\, \$v1999\, 
               \$v2007\, \$v1883\, \$258_len\, \$v1793\, \$278\, \$v1901\, 
               \$v1931\, \$328\, \$v1800\, \$v143\, \$277\, \$v1781\, \$295\, 
               \$333_i\, \$v128\, \$v1894\, \$260_i\, \$102_c\ : value(0 to 31) := (others => '0');
      variable \$arr1696_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1697_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1698_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1699_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1700_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1701_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1702_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1703_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1704_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v1873\); default_zero(\$102_c\); 
          default_zero(\$260_i\); default_zero(\$v1920\); 
          default_zero(\$v1641\); default_zero(\$v1965\); 
          default_zero(\$v1874\); default_zero(\$v1894\); 
          default_zero(\$v1907\); default_zero(\$v128\); 
          default_zero(\$268\); default_zero(\$333_i\); 
          default_zero(\$v2043\); default_zero(\$v1816\); 
          default_zero(\$v1806\); default_zero(\$v181\); 
          default_zero(\$295\); default_zero(\$v1720\); 
          default_zero(\$v1843\); default_zero(\$v106\); 
          default_zero(\$v2035\); default_zero(\$v1729\); 
          default_zero(\$v1781\); default_zero(\$277\); 
          default_zero(\$v1937\); default_zero(\$326\); 
          default_zero(\$v186\); default_zero(\$v143\); 
          default_zero(\$v1775\); default_zero(\$v1800\); 
          default_zero(\$v1737\); default_zero(\$v1783\); 
          default_zero(\$v1905\); default_zero(\$v130\); 
          default_zero(\$v1943\); default_zero(\$328\); 
          default_zero(\$v1931\); default_zero(\$v1979\); 
          default_zero(\$v2059\); default_zero(\$v2019\); 
          default_zero(\$v1901\); default_zero(\$278\); 
          default_zero(\$v2051\); default_zero(\$v1793\); 
          default_zero(\$258_len\); default_zero(\$v1970\); 
          default_zero(\$v104\); default_zero(\$v107\); 
          default_zero(\$v1821\); default_zero(\$v1711\); 
          default_zero(\$v1883\); default_zero(\$v1826\); 
          default_zero(\$v2007\); default_zero(\$v1999\); 
          default_zero(\$v1925\); default_zero(\$v1817\); 
          default_zero(\$269\); default_zero(\$v1838\); 
          default_zero(\$v1844\); default_zero(\$v1930\); 
          default_zero(\$74_i\); default_zero(\$v1893\); 
          default_zero(\$v1848\); default_zero(\$v1859\); 
          default_zero(\$v163\); default_zero(\$v1880\); 
          default_zero(\$v1749\); default_zero(\$v1878\); 
          default_zero(\$283\); default_zero(\$297\); default_zero(\$v145\); 
          default_zero(\$v170\); default_zero(\$265\); 
          default_zero(\$v1715\); default_zero(list_tail700_arg); 
          default_zero(\$v2067\); default_zero(\$v2015\); 
          default_zero(\$220_i\); default_zero(\$v1792\); 
          default_zero(\$v1782\); default_zero(\$v1993\); 
          default_zero(\$v1991\); default_zero(\$v147\); 
          default_zero(\$v1709\); default_zero(\$v158\); 
          default_zero(\$v1983\); default_zero(\$v1768\); 
          default_zero(\$v1935\); default_zero(\$v1994\); 
          default_zero(\$v116\); default_zero(\$v108\); 
          default_zero(\$v1911\); default_zero(\$v1854\); 
          default_zero(\$v115\); default_zero(\$v2014\); 
          default_zero(\$v1719\); default_zero(\$v1869\); 
          default_zero(\$292\); default_zero(\$v1951\); 
          default_zero(\$v148\); default_zero(\$v1741\); 
          default_zero(\$v185\); default_zero(\$264\); 
          default_zero(\$v1754\); default_zero(\$v1774\); 
          default_zero(\$v123\); default_zero(\$v1807\); 
          default_zero(aux7331672_arg); default_zero(\$v1756\); 
          default_zero(\$v1929\); default_zero(\$v1867\); 
          default_zero(\$v2055\); default_zero(\$v1788\); 
          default_zero(\$v1723\); default_zero(\$v1799\); 
          default_zero(\$v1727\); default_zero(\$v1940\); 
          default_zero(\$v184\); default_zero(\$v180\); 
          default_zero(\$v1795\); default_zero(\$327\); 
          default_zero(\$v110\); default_zero(\$v1891\); 
          default_zero(\$v1710\); default_zero(\$v1868\); 
          default_zero(\$v1853\); default_zero(aux7331672_result); 
          default_zero(\$v1956\); default_zero(\$v1881\); 
          default_zero(result1705); default_zero(\$v1898\); 
          default_zero(\$v1941\); default_zero(\$v1855\); 
          default_zero(\$v161\); default_zero(\$v2013\); 
          default_zero(get_int703_arg); default_zero(\$v1708\); 
          default_zero(\$v1753\); default_zero(loop3732_arg); 
          default_zero(\$89_i\); default_zero(\$324_c\); 
          default_zero(\$v1915\); default_zero(\$288_i\); 
          default_zero(\$267\); default_zero(\$v1955\); 
          default_zero(\$v2039\); default_zero(\$v1841\); 
          default_zero(\$71_x\); default_zero(\$v1808\); 
          default_zero(\$v129\); default_zero(\$222_i\); 
          default_zero(\$v1745\); default_zero(aux7331677_result); 
          default_zero(\$v198\); default_zero(\$v1899\); 
          default_zero(\$v1987\); default_zero(\$81_i\); 
          default_zero(\$v1975\); default_zero(\$v1822\); 
          default_zero(\$v2005\); default_zero(\$v1892\); 
          default_zero(\$v1969\); default_zero(\$325\); 
          default_zero(\$v1947\); default_zero(\$v2012\); 
          default_zero(\$v1971\); default_zero(\$v1879\); 
          default_zero(\$v1842\); default_zero(\$v1721\); 
          default_zero(\$v1887\); default_zero(\$v1728\); 
          default_zero(\$v1942\); default_zero(\$266\); 
          default_zero(\$v2047\); default_zero(\$v1830\); 
          default_zero(\$303\); default_zero(\$v1812\); 
          default_zero(\$v114\); default_zero(\$v1992\); 
          default_zero(\$v151\); default_zero(\$v1801\); 
          default_zero(\$v1863\); default_zero(\$v1760\); 
          default_zero(\$v1837\); default_zero(\$v179\); 
          default_zero(\$v105\); default_zero(\$v1840\); 
          default_zero(\$v1936\); default_zero(\$v113\); 
          default_zero(\$296\); default_zero(\$v146\); 
          default_zero(\$v1779\); default_zero(\$v2001\); 
          default_zero(\$v1802\); default_zero(\$v1794\); 
          default_zero(\$v1921\); default_zero(\$v1770\); 
          default_zero(\$v1733\); default_zero(\$v2027\); 
          default_zero(\$v1939\); default_zero(\$v2063\); 
          default_zero(\$v1852\); default_zero(\$v1839\); 
          default_zero(\$v111\); default_zero(\$v1900\); 
          default_zero(\$v1780\); default_zero(\$v1769\); 
          default_zero(\$v2023\); default_zero(\$v1998\); 
          default_zero(rdy1706); default_zero(\$v1906\); 
          default_zero(\$101_x\); default_zero(\$270_i\); 
          default_zero(\$v2031\); default_zero(\$286\); 
          default_zero(\$v1832\); default_zero(\$v2008\); 
          default_zero(\$274\); default_zero(\$v2000\); 
          default_zero(\$v1938\); default_zero(\$v112\); 
          default_zero(\$v125\); default_zero(\$279_i\); 
          default_zero(\$v1784\); default_zero(len); default_zero(\$v199\); 
          default_zero(\$v1831\); default_zero(\$99_x\); 
          default_zero(\$v124\); default_zero(\$v1722\); 
          default_zero(\$v1960\); default_zero(\$v1836\); 
          default_zero(\$v1764\); default_zero(\$v1916\); 
          default_zero(\$287\); default_zero(\$305_i\); 
          default_zero(\$76_x\); default_zero(\$v1755\); 
          default_zero(\$84_i\); default_zero(\$259_x\); 
          default_zero(\$87_i\); default_zero(aux7331677_arg); 
          default_zero(\$v2006\); default_zero(\$v1961\); 
          default_zero(\$v1882\); 
          rdy <= "1";
          rdy1706 := "0";
          \state\ <= compute1707;
          
        else if run = '1' then
          case \state\ is
          when \$234_forever7481664\ =>
            \state\ <= \$234_forever7481664\;
          when \$234_forever7481665\ =>
            \state\ <= \$234_forever7481665\;
          when \$234_forever7481666\ =>
            \state\ <= \$234_forever7481666\;
          when \$234_forever7481667\ =>
            \state\ <= \$234_forever7481667\;
          when \$234_forever7481668\ =>
            \state\ <= \$234_forever7481668\;
          when \$234_forever7481669\ =>
            \state\ <= \$234_forever7481669\;
          when \$234_forever7481670\ =>
            \state\ <= \$234_forever7481670\;
          when \$234_forever7481671\ =>
            \state\ <= \$234_forever7481671\;
          when \$234_forever7481673\ =>
            \state\ <= \$234_forever7481673\;
          when \$234_forever7481674\ =>
            \state\ <= \$234_forever7481674\;
          when \$234_forever7481675\ =>
            \state\ <= \$234_forever7481675\;
          when \$234_forever7481676\ =>
            \state\ <= \$234_forever7481676\;
          when \$310_forever7481665\ =>
            \state\ <= \$310_forever7481665\;
          when aux7331672 =>
            \$v1942\ := aux7331672_arg(72 to 107);
            \$v1943\ := \$v1942\(0 to 3);
            \$v1941\ := \$v1942\(4 to 35);
            case \$v1943\ is
            when "0001" =>
              \$v158\ := eclat_true;
              \$v1940\ := \$v158\;
              if \$v1940\(0) = '1' then
                \$v1938\ := aux7331672_arg(36 to 71);
                \$v1939\ := \$v1938\(0 to 3);
                \$v1930\ := \$v1938\(4 to 35);
                case \$v1939\ is
                when "0010" =>
                  \$81_i\ := \$v1930\(0 to 31);
                  \$v1936\ := "0010" & \$81_i\;
                  \$v1937\ := \$v1936\(0 to 3);
                  \$v1931\ := \$v1936\(4 to 35);
                  case \$v1937\ is
                  when "0010" =>
                    \$220_i\ := \$v1931\(0 to 31);
                    \$v1935\ := \$arr1697_ptr_take\;
                    if \$v1935\(0) = '1' then
                      \state\ <= q_wait1934;
                    else
                      \$arr1697_ptr_take\(0) := '1';
                      \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
                      \state\ <= pause_getI1932;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_rib expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$234_forever7481666\;
                  end case;
                when "0001" =>
                  aux7331672_result := eclat_add(aux7331672_arg(108 to 139) & "00000000000000000000000000000001");
                  len := aux7331672_result;
                  \$v1929\ := \$arr1700_ptr_take\;
                  if \$v1929\(0) = '1' then
                    \state\ <= q_wait1928;
                  else
                    \$arr1700_ptr_take\(0) := '1';
                    \$arr1700_ptr\ <= 0;
                    \state\ <= pause_getI1926;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("length"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$234_forever7481665\;
                end case;
              else
                aux7331672_result := aux7331672_arg(108 to 139);
                len := aux7331672_result;
                \$v1929\ := \$arr1700_ptr_take\;
                if \$v1929\(0) = '1' then
                  \state\ <= q_wait1928;
                else
                  \$arr1700_ptr_take\(0) := '1';
                  \$arr1700_ptr\ <= 0;
                  \state\ <= pause_getI1926;
                end if;
              end if;
            when others =>
              \$v158\ := eclat_false;
              \$v1940\ := \$v158\;
              if \$v1940\(0) = '1' then
                \$v1938\ := aux7331672_arg(36 to 71);
                \$v1939\ := \$v1938\(0 to 3);
                \$v1930\ := \$v1938\(4 to 35);
                case \$v1939\ is
                when "0010" =>
                  \$81_i\ := \$v1930\(0 to 31);
                  \$v1936\ := "0010" & \$81_i\;
                  \$v1937\ := \$v1936\(0 to 3);
                  \$v1931\ := \$v1936\(4 to 35);
                  case \$v1937\ is
                  when "0010" =>
                    \$220_i\ := \$v1931\(0 to 31);
                    \$v1935\ := \$arr1697_ptr_take\;
                    if \$v1935\(0) = '1' then
                      \state\ <= q_wait1934;
                    else
                      \$arr1697_ptr_take\(0) := '1';
                      \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
                      \state\ <= pause_getI1932;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_rib expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$234_forever7481666\;
                  end case;
                when "0001" =>
                  aux7331672_result := eclat_add(aux7331672_arg(108 to 139) & "00000000000000000000000000000001");
                  len := aux7331672_result;
                  \$v1929\ := \$arr1700_ptr_take\;
                  if \$v1929\(0) = '1' then
                    \state\ <= q_wait1928;
                  else
                    \$arr1700_ptr_take\(0) := '1';
                    \$arr1700_ptr\ <= 0;
                    \state\ <= pause_getI1926;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("length"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$234_forever7481665\;
                end case;
              else
                aux7331672_result := aux7331672_arg(108 to 139);
                len := aux7331672_result;
                \$v1929\ := \$arr1700_ptr_take\;
                if \$v1929\(0) = '1' then
                  \state\ <= q_wait1928;
                else
                  \$arr1700_ptr_take\(0) := '1';
                  \$arr1700_ptr\ <= 0;
                  \state\ <= pause_getI1926;
                end if;
              end if;
            end case;
          when aux7331677 =>
            \$v1843\ := aux7331677_arg(72 to 107);
            \$v1844\ := \$v1843\(0 to 3);
            \$v1842\ := \$v1843\(4 to 35);
            case \$v1844\ is
            when "0001" =>
              \$303\ := eclat_true;
              \$v1841\ := \$303\;
              if \$v1841\(0) = '1' then
                \$v1839\ := aux7331677_arg(36 to 71);
                \$v1840\ := \$v1839\(0 to 3);
                \$v1831\ := \$v1839\(4 to 35);
                case \$v1840\ is
                when "0010" =>
                  \$305_i\ := \$v1831\(0 to 31);
                  \$v1837\ := "0010" & \$305_i\;
                  \$v1838\ := \$v1837\(0 to 3);
                  \$v1832\ := \$v1837\(4 to 35);
                  case \$v1838\ is
                  when "0010" =>
                    \$220_i\ := \$v1832\(0 to 31);
                    \$v1836\ := \$arr1697_ptr_take\;
                    if \$v1836\(0) = '1' then
                      \state\ <= q_wait1835;
                    else
                      \$arr1697_ptr_take\(0) := '1';
                      \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
                      \state\ <= pause_getI1833;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_rib expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$234_forever7481666\;
                  end case;
                when "0001" =>
                  aux7331677_result := eclat_add(aux7331677_arg(108 to 139) & "00000000000000000000000000000001");
                  \$258_len\ := aux7331677_result;
                  \$v1830\ := \$arr1700_ptr_take\;
                  if \$v1830\(0) = '1' then
                    \state\ <= q_wait1829;
                  else
                    \$arr1700_ptr_take\(0) := '1';
                    \$arr1700_ptr\ <= 0;
                    \state\ <= pause_getI1827;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("length"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$310_forever7481665\;
                end case;
              else
                aux7331677_result := aux7331677_arg(108 to 139);
                \$258_len\ := aux7331677_result;
                \$v1830\ := \$arr1700_ptr_take\;
                if \$v1830\(0) = '1' then
                  \state\ <= q_wait1829;
                else
                  \$arr1700_ptr_take\(0) := '1';
                  \$arr1700_ptr\ <= 0;
                  \state\ <= pause_getI1827;
                end if;
              end if;
            when others =>
              \$303\ := eclat_false;
              \$v1841\ := \$303\;
              if \$v1841\(0) = '1' then
                \$v1839\ := aux7331677_arg(36 to 71);
                \$v1840\ := \$v1839\(0 to 3);
                \$v1831\ := \$v1839\(4 to 35);
                case \$v1840\ is
                when "0010" =>
                  \$305_i\ := \$v1831\(0 to 31);
                  \$v1837\ := "0010" & \$305_i\;
                  \$v1838\ := \$v1837\(0 to 3);
                  \$v1832\ := \$v1837\(4 to 35);
                  case \$v1838\ is
                  when "0010" =>
                    \$220_i\ := \$v1832\(0 to 31);
                    \$v1836\ := \$arr1697_ptr_take\;
                    if \$v1836\(0) = '1' then
                      \state\ <= q_wait1835;
                    else
                      \$arr1697_ptr_take\(0) := '1';
                      \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
                      \state\ <= pause_getI1833;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_rib expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$234_forever7481666\;
                  end case;
                when "0001" =>
                  aux7331677_result := eclat_add(aux7331677_arg(108 to 139) & "00000000000000000000000000000001");
                  \$258_len\ := aux7331677_result;
                  \$v1830\ := \$arr1700_ptr_take\;
                  if \$v1830\(0) = '1' then
                    \state\ <= q_wait1829;
                  else
                    \$arr1700_ptr_take\(0) := '1';
                    \$arr1700_ptr\ <= 0;
                    \state\ <= pause_getI1827;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("length"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$310_forever7481665\;
                end case;
              else
                aux7331677_result := aux7331677_arg(108 to 139);
                \$258_len\ := aux7331677_result;
                \$v1830\ := \$arr1700_ptr_take\;
                if \$v1830\(0) = '1' then
                  \state\ <= q_wait1829;
                else
                  \$arr1700_ptr_take\(0) := '1';
                  \$arr1700_ptr\ <= 0;
                  \state\ <= pause_getI1827;
                end if;
              end if;
            end case;
          when get_int703 =>
            \$v1745\ := \$arr1702_ptr_take\;
            if \$v1745\(0) = '1' then
              \state\ <= q_wait1744;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1742;
            end if;
          when list_tail700 =>
            \$v1728\ := eclat_eq("00000000000000000000000000000000" & list_tail700_arg(32 to 63));
            if \$v1728\(0) = '1' then
              \$v1708\ := list_tail700_arg(0 to 31);
              
              \state\ <= list_tail700;
            else
              \$v1727\ := \$arr1697_ptr_take\;
              if \$v1727\(0) = '1' then
                \state\ <= q_wait1726;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
                \state\ <= pause_getI1724;
              end if;
            end if;
          when loop3732 =>
            \$v1987\ := \$arr1702_ptr_take\;
            if \$v1987\(0) = '1' then
              \state\ <= q_wait1986;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1984;
            end if;
          when pause_getI1712 =>
            \state\ <= pause_getII1713;
          when pause_getI1716 =>
            \state\ <= pause_getII1717;
          when pause_getI1724 =>
            \state\ <= pause_getII1725;
          when pause_getI1734 =>
            \state\ <= pause_getII1735;
          when pause_getI1738 =>
            \state\ <= pause_getII1739;
          when pause_getI1742 =>
            \state\ <= pause_getII1743;
          when pause_getI1746 =>
            \state\ <= pause_getII1747;
          when pause_getI1771 =>
            \state\ <= pause_getII1772;
          when pause_getI1776 =>
            \state\ <= pause_getII1777;
          when pause_getI1785 =>
            \state\ <= pause_getII1786;
          when pause_getI1789 =>
            \state\ <= pause_getII1790;
          when pause_getI1809 =>
            \state\ <= pause_getII1810;
          when pause_getI1813 =>
            \state\ <= pause_getII1814;
          when pause_getI1823 =>
            \state\ <= pause_getII1824;
          when pause_getI1827 =>
            \state\ <= pause_getII1828;
          when pause_getI1833 =>
            \state\ <= pause_getII1834;
          when pause_getI1845 =>
            \state\ <= pause_getII1846;
          when pause_getI1870 =>
            \state\ <= pause_getII1871;
          when pause_getI1875 =>
            \state\ <= pause_getII1876;
          when pause_getI1884 =>
            \state\ <= pause_getII1885;
          when pause_getI1888 =>
            \state\ <= pause_getII1889;
          when pause_getI1908 =>
            \state\ <= pause_getII1909;
          when pause_getI1912 =>
            \state\ <= pause_getII1913;
          when pause_getI1922 =>
            \state\ <= pause_getII1923;
          when pause_getI1926 =>
            \state\ <= pause_getII1927;
          when pause_getI1932 =>
            \state\ <= pause_getII1933;
          when pause_getI1944 =>
            \state\ <= pause_getII1945;
          when pause_getI1948 =>
            \state\ <= pause_getII1949;
          when pause_getI1962 =>
            \state\ <= pause_getII1963;
          when pause_getI1966 =>
            \state\ <= pause_getII1967;
          when pause_getI1976 =>
            \state\ <= pause_getII1977;
          when pause_getI1980 =>
            \state\ <= pause_getII1981;
          when pause_getI1984 =>
            \state\ <= pause_getII1985;
          when pause_getII1713 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1641\ := \$arr1697_value\;
            \$v1710\ := \$v1641\(36 to 71);
            \$v1711\ := \$v1710\(0 to 3);
            \$v1709\ := \$v1710\(4 to 35);
            case \$v1711\ is
            when "0010" =>
              \$333_i\ := \$v1709\(0 to 31);
              \$v108\ := \$333_i\;
              \$v110\ := \$v108\ & eclat_sub(list_tail700_arg(32 to 63) & "00000000000000000000000000000001");
              list_tail700_arg := \$v110\;
              \state\ <= list_tail700;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481664\;
            end case;
          when pause_getII1717 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v107\ := \$arr1697_value\;
            \state\ <= list_tail700;
          when pause_getII1725 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v104\ := \$arr1697_value\;
            \$v105\ := \$v104\(36 to 71);
            \$v1722\ := \$v105\;
            \$v1723\ := \$v1722\(0 to 3);
            \$v1721\ := \$v1722\(4 to 35);
            case \$v1723\ is
            when "0010" =>
              \$v106\ := eclat_true;
              \$v1720\ := \$v106\;
              if \$v1720\(0) = '1' then
                \$v1715\ := \$arr1697_ptr_take\;
                if \$v1715\(0) = '1' then
                  \state\ <= q_wait1714;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
                  \state\ <= pause_getI1712;
                end if;
              else
                \$v1719\ := \$arr1697_ptr_take\;
                if \$v1719\(0) = '1' then
                  \state\ <= q_wait1718;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
                  \state\ <= pause_getI1716;
                end if;
              end if;
            when others =>
              \$v106\ := eclat_false;
              \$v1720\ := \$v106\;
              if \$v1720\(0) = '1' then
                \$v1715\ := \$arr1697_ptr_take\;
                if \$v1715\(0) = '1' then
                  \state\ <= q_wait1714;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
                  \state\ <= pause_getI1712;
                end if;
              else
                \$v1719\ := \$arr1697_ptr_take\;
                if \$v1719\(0) = '1' then
                  \state\ <= q_wait1718;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
                  \state\ <= pause_getI1716;
                end if;
              end if;
            end case;
          when pause_getII1735 =>
            \$arr1702_ptr_take\(0) := '0';
            \$327\ := \$arr1702_value\;
            \$326\ := \$327\ & "00000000000000000000000000000001";
            \$325\ := eclat_add(\$326\);
            \$v1733\ := \$arr1702_ptr_take\;
            if \$v1733\(0) = '1' then
              \state\ <= q_wait1732;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= \$325\;
              \state\ <= pause_setI1730;
            end if;
          when pause_getII1739 =>
            \$arr1696_ptr_take\(0) := '0';
            \$324_c\ := \$arr1696_value\;
            \$v1737\ := \$arr1702_ptr_take\;
            if \$v1737\(0) = '1' then
              \state\ <= q_wait1736;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1734;
            end if;
          when pause_getII1743 =>
            \$arr1702_ptr_take\(0) := '0';
            \$328\ := \$arr1702_value\;
            \$v1741\ := \$arr1696_ptr_take\;
            if \$v1741\(0) = '1' then
              \state\ <= q_wait1740;
            else
              \$arr1696_ptr_take\(0) := '1';
              \$arr1696_ptr\ <= to_integer(unsigned(\$328\));
              \state\ <= pause_getI1738;
            end if;
          when pause_getII1747 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v199\ := \$arr1700_value\;
            loop3732_arg := \$v199\;
            \state\ <= loop3732;
          when pause_getII1772 =>
            \$arr1701_ptr_take\(0) := '0';
            \$267\ := \$arr1701_value\;
            \$266\ := "0010" & \$267\;
            \$v1769\ := eclat_add(\$259_x\ & "00000000000000000000000000000010");
            \$v1770\ := "00000000000000000000000000000000";
            \$265\ := "0010" & \$v1769\ & \$266\ & "0001" & \$v1770\;
            \$v1768\ := \$arr1697_ptr_take\;
            if \$v1768\(0) = '1' then
              \state\ <= q_wait1767;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$260_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= \$265\;
              \state\ <= pause_setI1765;
            end if;
          when pause_getII1777 =>
            \$arr1701_ptr_take\(0) := '0';
            \$269\ := \$arr1701_value\;
            \$268\ := \$269\ & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
            \$264\ := eclat_eq(\$268\);
            \$v1775\ := \$264\;
            if \$v1775\(0) = '1' then
              \$v1760\ := \$arr1697_ptr_take\;
              if \$v1760\(0) = '1' then
                \state\ <= q_wait1759;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$v1754\ := eclat_add(\$259_x\ & "00000000000000000000000000000010");
                \$v1755\ := "00000000000000000000000000000000";
                \$v1756\ := "00000000000000000000000000000000";
                \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$260_i\ & "00000000000000000000000000000001")));
                \$arr1697_write_request\ <= '1';
                \$arr1697_write\ <= "0010" & \$v1754\ & "0001" & \$v1755\ & "0001" & \$v1756\;
                \state\ <= pause_setI1757;
              end if;
            else
              \$v1774\ := \$arr1701_ptr_take\;
              if \$v1774\(0) = '1' then
                \state\ <= q_wait1773;
              else
                \$arr1701_ptr_take\(0) := '1';
                \$arr1701_ptr\ <= 0;
                \state\ <= pause_getI1771;
              end if;
            end if;
          when pause_getII1786 =>
            \$arr1701_ptr_take\(0) := '0';
            \$278\ := \$arr1701_value\;
            \$274\ := \$277\ & \$278\;
            \$259_x\ := eclat_if(eclat_gt(\$274\(32 to 63) & \$274\(0 to 31)) & \$274\(32 to 63) & \$274\(0 to 31));
            \$v1784\ := eclat_add(\$259_x\ & "00000000000000000000000000000010");
            \$v1782\ := "0010" & \$v1784\;
            \$v1783\ := \$v1782\(0 to 3);
            \$v1781\ := \$v1782\(4 to 35);
            case \$v1783\ is
            when "0010" =>
              \$270_i\ := \$v1781\(0 to 31);
              \$260_i\ := \$270_i\;
              \$v1780\ := eclat_lt(\$260_i\ & eclat_sub(eclat_div(X"0000" & X"2328" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1780\(0) = '1' then
                \$v1779\ := \$arr1701_ptr_take\;
                if \$v1779\(0) = '1' then
                  \state\ <= q_wait1778;
                else
                  \$arr1701_ptr_take\(0) := '1';
                  \$arr1701_ptr\ <= 0;
                  \state\ <= pause_getI1776;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow push_word_stbl "));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$234_forever7481673\;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481674\;
            end case;
          when pause_getII1790 =>
            \$arr1700_ptr_take\(0) := '0';
            \$277\ := \$arr1700_value\;
            \$v1788\ := \$arr1701_ptr_take\;
            if \$v1788\(0) = '1' then
              \state\ <= q_wait1787;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1785;
            end if;
          when pause_getII1810 =>
            \$arr1701_ptr_take\(0) := '0';
            \$287\ := \$arr1701_value\;
            \$283\ := \$286\ & \$287\;
            \$279_i\ := eclat_if(eclat_gt(\$283\(32 to 63) & \$283\(0 to 31)) & \$283\(32 to 63) & \$283\(0 to 31));
            \$v1808\ := eclat_lt(\$279_i\ & eclat_sub(eclat_div(X"0000" & X"2328" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
            if \$v1808\(0) = '1' then
              \$v1807\ := eclat_eq(\$279_i\ & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001"));
              if \$v1807\(0) = '1' then
                \$v1799\ := \$arr1697_ptr_take\;
                if \$v1799\(0) = '1' then
                  \state\ <= q_wait1798;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$v1793\ := "00000000000000000000000000000011";
                  \$v1794\ := "00000000000000000000000000000000";
                  \$v1795\ := "00000000000000000000000000000010";
                  \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$279_i\ & "00000000000000000000000000000010")));
                  \$arr1697_write_request\ <= '1';
                  \$arr1697_write\ <= "0010" & \$v1793\ & "0001" & \$v1794\ & "0001" & \$v1795\;
                  \state\ <= pause_setI1796;
                end if;
              else
                \$v1806\ := \$arr1697_ptr_take\;
                if \$v1806\(0) = '1' then
                  \state\ <= q_wait1805;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$v1800\ := "00000000000000000000000000000011";
                  \$v1801\ := eclat_add(\$279_i\ & "00000000000000000000000000000001");
                  \$v1802\ := "00000000000000000000000000000010";
                  \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$279_i\ & "00000000000000000000000000000010")));
                  \$arr1697_write_request\ <= '1';
                  \$arr1697_write\ <= "0010" & \$v1800\ & "0010" & \$v1801\ & "0001" & \$v1802\;
                  \state\ <= pause_setI1803;
                end if;
              end if;
            else
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("stack overflow push2_symtbl_word"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481675\;
            end if;
          when pause_getII1814 =>
            \$arr1700_ptr_take\(0) := '0';
            \$286\ := \$arr1700_value\;
            \$v1812\ := \$arr1701_ptr_take\;
            if \$v1812\(0) = '1' then
              \state\ <= q_wait1811;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1809;
            end if;
          when pause_getII1824 =>
            \$arr1701_ptr_take\(0) := '0';
            \$296\ := \$arr1701_value\;
            \$292\ := \$295\ & \$296\;
            \$288_i\ := eclat_if(eclat_gt(\$292\(32 to 63) & \$292\(0 to 31)) & \$292\(32 to 63) & \$292\(0 to 31));
            \$v1822\ := eclat_lt(\$288_i\ & X"0000" & X"2328");
            if \$v1822\(0) = '1' then
              \$v1821\ := \$arr1697_ptr_take\;
              if \$v1821\(0) = '1' then
                \state\ <= q_wait1820;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$v1817\ := "00000000000000000000000000000011";
                \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$288_i\ & "00000000000000000000000000000001")));
                \$arr1697_write_request\ <= '1';
                \$arr1697_write\ <= "0010" & loop3732_arg & "0001" & \$258_len\ & "0001" & \$v1817\;
                \state\ <= pause_setI1818;
              end if;
            else
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("stack overflow push_symtbl_rib"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481676\;
            end if;
          when pause_getII1828 =>
            \$arr1700_ptr_take\(0) := '0';
            \$295\ := \$arr1700_value\;
            \$v1826\ := \$arr1701_ptr_take\;
            if \$v1826\(0) = '1' then
              \state\ <= q_wait1825;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1823;
            end if;
          when pause_getII1834 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v161\ := \$arr1697_value\;
            \$v163\ := \$v161\ & eclat_add(aux7331677_arg(108 to 139) & "00000000000000000000000000000001");
            aux7331677_arg := \$v163\;
            \state\ <= aux7331677;
          when pause_getII1846 =>
            \$arr1697_ptr_take\(0) := '0';
            \$297\ := \$arr1697_value\;
            aux7331677_arg := \$297\ & "00000000000000000000000000000000";
            \state\ <= aux7331677;
          when pause_getII1871 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v147\ := \$arr1701_value\;
            \$v148\ := "0010" & \$v147\;
            \$v1868\ := eclat_add(\$76_x\ & "00000000000000000000000000000010");
            \$v1869\ := "00000000000000000000000000000000";
            \$v151\ := "0010" & \$v1868\ & \$v148\ & "0001" & \$v1869\;
            \$v1867\ := \$arr1697_ptr_take\;
            if \$v1867\(0) = '1' then
              \state\ <= q_wait1866;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$84_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= \$v151\;
              \state\ <= pause_setI1864;
            end if;
          when pause_getII1876 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v143\ := \$arr1701_value\;
            \$v145\ := \$v143\ & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
            \$v146\ := eclat_eq(\$v145\);
            \$v1874\ := \$v146\;
            if \$v1874\(0) = '1' then
              \$v1859\ := \$arr1697_ptr_take\;
              if \$v1859\(0) = '1' then
                \state\ <= q_wait1858;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$v1853\ := eclat_add(\$76_x\ & "00000000000000000000000000000010");
                \$v1854\ := "00000000000000000000000000000000";
                \$v1855\ := "00000000000000000000000000000000";
                \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$84_i\ & "00000000000000000000000000000001")));
                \$arr1697_write_request\ <= '1';
                \$arr1697_write\ <= "0010" & \$v1853\ & "0001" & \$v1854\ & "0001" & \$v1855\;
                \state\ <= pause_setI1856;
              end if;
            else
              \$v1873\ := \$arr1701_ptr_take\;
              if \$v1873\(0) = '1' then
                \state\ <= q_wait1872;
              else
                \$arr1701_ptr_take\(0) := '1';
                \$arr1701_ptr\ <= 0;
                \state\ <= pause_getI1870;
              end if;
            end if;
          when pause_getII1885 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v180\ := \$arr1701_value\;
            \$v181\ := \$v179\ & \$v180\;
            \$76_x\ := eclat_if(eclat_gt(\$v181\(32 to 63) & \$v181\(0 to 31)) & \$v181\(32 to 63) & \$v181\(0 to 31));
            \$v1883\ := eclat_add(\$76_x\ & "00000000000000000000000000000010");
            \$v1881\ := "0010" & \$v1883\;
            \$v1882\ := \$v1881\(0 to 3);
            \$v1880\ := \$v1881\(4 to 35);
            case \$v1882\ is
            when "0010" =>
              \$222_i\ := \$v1880\(0 to 31);
              \$84_i\ := \$222_i\;
              \$v1879\ := eclat_lt(\$84_i\ & eclat_sub(eclat_div(X"0000" & X"2328" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1879\(0) = '1' then
                \$v1878\ := \$arr1701_ptr_take\;
                if \$v1878\(0) = '1' then
                  \state\ <= q_wait1877;
                else
                  \$arr1701_ptr_take\(0) := '1';
                  \$arr1701_ptr\ <= 0;
                  \state\ <= pause_getI1875;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow push_word_stbl "));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$234_forever7481668\;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481669\;
            end case;
          when pause_getII1889 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v179\ := \$arr1700_value\;
            \$v1887\ := \$arr1701_ptr_take\;
            if \$v1887\(0) = '1' then
              \state\ <= q_wait1886;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1884;
            end if;
          when pause_getII1909 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v129\ := \$arr1701_value\;
            \$v130\ := \$v128\ & \$v129\;
            \$87_i\ := eclat_if(eclat_gt(\$v130\(32 to 63) & \$v130\(0 to 31)) & \$v130\(32 to 63) & \$v130\(0 to 31));
            \$v1907\ := eclat_lt(\$87_i\ & eclat_sub(eclat_div(X"0000" & X"2328" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
            if \$v1907\(0) = '1' then
              \$v1906\ := eclat_eq(\$87_i\ & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001"));
              if \$v1906\(0) = '1' then
                \$v1898\ := \$arr1697_ptr_take\;
                if \$v1898\(0) = '1' then
                  \state\ <= q_wait1897;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$v1892\ := "00000000000000000000000000000011";
                  \$v1893\ := "00000000000000000000000000000000";
                  \$v1894\ := "00000000000000000000000000000010";
                  \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$87_i\ & "00000000000000000000000000000010")));
                  \$arr1697_write_request\ <= '1';
                  \$arr1697_write\ <= "0010" & \$v1892\ & "0001" & \$v1893\ & "0001" & \$v1894\;
                  \state\ <= pause_setI1895;
                end if;
              else
                \$v1905\ := \$arr1697_ptr_take\;
                if \$v1905\(0) = '1' then
                  \state\ <= q_wait1904;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$v1899\ := "00000000000000000000000000000011";
                  \$v1900\ := eclat_add(\$87_i\ & "00000000000000000000000000000001");
                  \$v1901\ := "00000000000000000000000000000010";
                  \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$87_i\ & "00000000000000000000000000000010")));
                  \$arr1697_write_request\ <= '1';
                  \$arr1697_write\ <= "0010" & \$v1899\ & "0010" & \$v1900\ & "0001" & \$v1901\;
                  \state\ <= pause_setI1902;
                end if;
              end if;
            else
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("stack overflow push2_symtbl_word"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481670\;
            end if;
          when pause_getII1913 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v128\ := \$arr1700_value\;
            \$v1911\ := \$arr1701_ptr_take\;
            if \$v1911\(0) = '1' then
              \state\ <= q_wait1910;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1908;
            end if;
          when pause_getII1923 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v124\ := \$arr1701_value\;
            \$v125\ := \$v123\ & \$v124\;
            \$89_i\ := eclat_if(eclat_gt(\$v125\(32 to 63) & \$v125\(0 to 31)) & \$v125\(32 to 63) & \$v125\(0 to 31));
            \$v1921\ := eclat_lt(\$89_i\ & X"0000" & X"2328");
            if \$v1921\(0) = '1' then
              \$v1920\ := \$arr1697_ptr_take\;
              if \$v1920\(0) = '1' then
                \state\ <= q_wait1919;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$v1916\ := "00000000000000000000000000000011";
                \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$89_i\ & "00000000000000000000000000000001")));
                \$arr1697_write_request\ <= '1';
                \$arr1697_write\ <= "0010" & loop3732_arg & "0001" & len & "0001" & \$v1916\;
                \state\ <= pause_setI1917;
              end if;
            else
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("stack overflow push_symtbl_rib"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481671\;
            end if;
          when pause_getII1927 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v123\ := \$arr1700_value\;
            \$v1925\ := \$arr1701_ptr_take\;
            if \$v1925\(0) = '1' then
              \state\ <= q_wait1924;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1922;
            end if;
          when pause_getII1933 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v161\ := \$arr1697_value\;
            \$v163\ := \$v161\ & eclat_add(aux7331672_arg(108 to 139) & "00000000000000000000000000000001");
            aux7331672_arg := \$v163\;
            \state\ <= aux7331672;
          when pause_getII1945 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v170\ := \$arr1697_value\;
            aux7331672_arg := \$v170\ & "00000000000000000000000000000000";
            \state\ <= aux7331672;
          when pause_getII1949 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v198\ := \$arr1700_value\;
            loop3732_arg := \$v198\;
            \state\ <= loop3732;
          when pause_getII1963 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v185\ := \$arr1700_value\;
            \$v186\ := \$v184\ & \$v185\;
            \$74_i\ := eclat_if(eclat_gt(\$v186\(32 to 63) & \$v186\(0 to 31)) & \$v186\(32 to 63) & \$v186\(0 to 31));
            \$v1961\ := eclat_lt(\$74_i\ & eclat_sub(eclat_div(X"0000" & X"2328" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
            if \$v1961\(0) = '1' then
              \$v1960\ := \$arr1697_ptr_take\;
              if \$v1960\(0) = '1' then
                \state\ <= q_wait1959;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$v1956\ := "00000000000000000000000000000000";
                \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$74_i\ & "00000000000000000000000000000001")));
                \$arr1697_write_request\ <= '1';
                \$arr1697_write\ <= "0001" & \$71_x\ & "0010" & loop3732_arg & "0001" & \$v1956\;
                \state\ <= pause_setI1957;
              end if;
            else
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("stack overflow push_symtbl_word_accum"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$234_forever7481667\;
            end if;
          when pause_getII1967 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v184\ := \$arr1701_value\;
            \$v1965\ := \$arr1700_ptr_take\;
            if \$v1965\(0) = '1' then
              \state\ <= q_wait1964;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1962;
            end if;
          when pause_getII1977 =>
            \$arr1702_ptr_take\(0) := '0';
            \$v112\ := \$arr1702_value\;
            \$v113\ := \$v112\ & "00000000000000000000000000000001";
            \$v114\ := eclat_add(\$v113\);
            \$v1975\ := \$arr1702_ptr_take\;
            if \$v1975\(0) = '1' then
              \state\ <= q_wait1974;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= \$v114\;
              \state\ <= pause_setI1972;
            end if;
          when pause_getII1981 =>
            \$arr1696_ptr_take\(0) := '0';
            \$102_c\ := \$arr1696_value\;
            \$v1979\ := \$arr1702_ptr_take\;
            if \$v1979\(0) = '1' then
              \state\ <= q_wait1978;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1976;
            end if;
          when pause_getII1985 =>
            \$arr1702_ptr_take\(0) := '0';
            \$v111\ := \$arr1702_value\;
            \$v1983\ := \$arr1696_ptr_take\;
            if \$v1983\(0) = '1' then
              \state\ <= q_wait1982;
            else
              \$arr1696_ptr_take\(0) := '1';
              \$arr1696_ptr\ <= to_integer(unsigned(\$v111\));
              \state\ <= pause_getI1980;
            end if;
          when pause_setI1730 =>
            \$arr1702_write_request\ <= '0';
            \state\ <= pause_setII1731;
          when pause_setI1750 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII1751;
          when pause_setI1757 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1758;
          when pause_setI1761 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII1762;
          when pause_setI1765 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1766;
          when pause_setI1796 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1797;
          when pause_setI1803 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1804;
          when pause_setI1818 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1819;
          when pause_setI1849 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII1850;
          when pause_setI1856 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1857;
          when pause_setI1860 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII1861;
          when pause_setI1864 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1865;
          when pause_setI1895 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1896;
          when pause_setI1902 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1903;
          when pause_setI1917 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1918;
          when pause_setI1952 =>
            \$arr1700_write_request\ <= '0';
            \state\ <= pause_setII1953;
          when pause_setI1957 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1958;
          when pause_setI1972 =>
            \$arr1702_write_request\ <= '0';
            \state\ <= pause_setII1973;
          when pause_setI1988 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII1989;
          when pause_setI1995 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII1996;
          when pause_setI2002 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII2003;
          when pause_setI2009 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII2010;
          when pause_setI2016 =>
            \$arr1697_write_request\ <= '0';
            \state\ <= pause_setII2017;
          when pause_setI2020 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2021;
          when pause_setI2024 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2025;
          when pause_setI2028 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2029;
          when pause_setI2032 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2033;
          when pause_setI2036 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2037;
          when pause_setI2040 =>
            \$arr1704_write_request\ <= '0';
            \state\ <= pause_setII2041;
          when pause_setI2044 =>
            \$arr1703_write_request\ <= '0';
            \state\ <= pause_setII2045;
          when pause_setI2048 =>
            \$arr1702_write_request\ <= '0';
            \state\ <= pause_setII2049;
          when pause_setI2052 =>
            \$arr1701_write_request\ <= '0';
            \state\ <= pause_setII2053;
          when pause_setI2056 =>
            \$arr1700_write_request\ <= '0';
            \state\ <= pause_setII2057;
          when pause_setI2060 =>
            \$arr1699_write_request\ <= '0';
            \state\ <= pause_setII2061;
          when pause_setI2064 =>
            \$arr1698_write_request\ <= '0';
            \state\ <= pause_setII2065;
          when pause_setII1731 =>
            \$arr1702_ptr_take\(0) := '0';
            \$v115\ := \$324_c\;
            \$v116\ := \$v115\ & X"000000" & X"23";
            \$101_x\ := eclat_sub(\$v116\);
            \$99_x\ := eclat_if(eclat_lt(\$101_x\ & "00000000000000000000000000000000") & X"000000" & X"39" & \$101_x\);
            \$v1729\ := eclat_lt(\$99_x\ & X"000000" & X"2e");
            if \$v1729\(0) = '1' then
              \state\ <= get_int703;
            else
              get_int703_arg := eclat_sub(eclat_add(eclat_mult(get_int703_arg & X"000000" & X"2e") & \$99_x\) & X"000000" & X"2e");
              \state\ <= get_int703;
            end if;
          when pause_setII1751 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v1749\ := \$arr1700_ptr_take\;
            if \$v1749\(0) = '1' then
              \state\ <= q_wait1748;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1746;
            end if;
          when pause_setII1758 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1753\ := \$arr1701_ptr_take\;
            if \$v1753\(0) = '1' then
              \state\ <= q_wait1752;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$260_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1750;
            end if;
          when pause_setII1762 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v1749\ := \$arr1700_ptr_take\;
            if \$v1749\(0) = '1' then
              \state\ <= q_wait1748;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1746;
            end if;
          when pause_setII1766 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1764\ := \$arr1701_ptr_take\;
            if \$v1764\(0) = '1' then
              \state\ <= q_wait1763;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$260_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1761;
            end if;
          when pause_setII1797 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1792\ := \$arr1700_ptr_take\;
            if \$v1792\(0) = '1' then
              \state\ <= q_wait1791;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1789;
            end if;
          when pause_setII1804 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1792\ := \$arr1700_ptr_take\;
            if \$v1792\(0) = '1' then
              \state\ <= q_wait1791;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1789;
            end if;
          when pause_setII1819 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1816\ := \$arr1700_ptr_take\;
            if \$v1816\(0) = '1' then
              \state\ <= q_wait1815;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1813;
            end if;
          when pause_setII1850 =>
            \$arr1701_ptr_take\(0) := '0';
            \state\ <= loop3732;
          when pause_setII1857 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1852\ := \$arr1701_ptr_take\;
            if \$v1852\(0) = '1' then
              \state\ <= q_wait1851;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$84_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1849;
            end if;
          when pause_setII1861 =>
            \$arr1701_ptr_take\(0) := '0';
            \state\ <= loop3732;
          when pause_setII1865 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1863\ := \$arr1701_ptr_take\;
            if \$v1863\(0) = '1' then
              \state\ <= q_wait1862;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$84_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1860;
            end if;
          when pause_setII1896 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1891\ := \$arr1700_ptr_take\;
            if \$v1891\(0) = '1' then
              \state\ <= q_wait1890;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1888;
            end if;
          when pause_setII1903 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1891\ := \$arr1700_ptr_take\;
            if \$v1891\(0) = '1' then
              \state\ <= q_wait1890;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1888;
            end if;
          when pause_setII1918 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1915\ := \$arr1700_ptr_take\;
            if \$v1915\(0) = '1' then
              \state\ <= q_wait1914;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1912;
            end if;
          when pause_setII1953 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v1951\ := \$arr1700_ptr_take\;
            if \$v1951\(0) = '1' then
              \state\ <= q_wait1950;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1948;
            end if;
          when pause_setII1958 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1955\ := \$arr1700_ptr_take\;
            if \$v1955\(0) = '1' then
              \state\ <= q_wait1954;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr_write\ <= 0;
              \$arr1700_write_request\ <= '1';
              \$arr1700_write\ <= eclat_add(\$74_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1952;
            end if;
          when pause_setII1973 =>
            \$arr1702_ptr_take\(0) := '0';
            \$71_x\ := \$102_c\;
            \$v1971\ := eclat_eq(\$71_x\ & X"000000" & X"2c");
            if \$v1971\(0) = '1' then
              \$v1848\ := \$arr1697_ptr_take\;
              if \$v1848\(0) = '1' then
                \state\ <= q_wait1847;
              else
                \$arr1697_ptr_take\(0) := '1';
                \$arr1697_ptr\ <= to_integer(unsigned(loop3732_arg));
                \state\ <= pause_getI1845;
              end if;
            else
              \$v1970\ := eclat_eq(\$71_x\ & X"000000" & X"3b");
              if \$v1970\(0) = '1' then
                \$v1947\ := \$arr1697_ptr_take\;
                if \$v1947\(0) = '1' then
                  \state\ <= q_wait1946;
                else
                  \$arr1697_ptr_take\(0) := '1';
                  \$arr1697_ptr\ <= to_integer(unsigned(loop3732_arg));
                  \state\ <= pause_getI1944;
                end if;
              else
                \$v1969\ := \$arr1701_ptr_take\;
                if \$v1969\(0) = '1' then
                  \state\ <= q_wait1968;
                else
                  \$arr1701_ptr_take\(0) := '1';
                  \$arr1701_ptr\ <= 0;
                  \state\ <= pause_getI1966;
                end if;
              end if;
            end if;
          when pause_setII1989 =>
            \$arr1701_ptr_take\(0) := '0';
            result1705 := eclat_unit;
            eclat_print_string(of_string("Test"));
            
            rdy1706 := eclat_true;
            \state\ <= compute1707;
          when pause_setII1996 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1991\ := \$arr1701_ptr_take\;
            if \$v1991\(0) = '1' then
              \state\ <= q_wait1990;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= "00000000000000000000000000000011";
              \state\ <= pause_setI1988;
            end if;
          when pause_setII2003 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v1998\ := \$arr1697_ptr_take\;
            if \$v1998\(0) = '1' then
              \state\ <= q_wait1997;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1992\ := "00000000000000000000000000000001";
              \$v1993\ := "00000000000000000000000000000010";
              \$v1994\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 3;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1992\ & "0010" & \$v1993\ & "0001" & \$v1994\;
              \state\ <= pause_setI1995;
            end if;
          when pause_setII2010 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v2005\ := \$arr1697_ptr_take\;
            if \$v2005\(0) = '1' then
              \state\ <= q_wait2004;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1999\ := "00000000000000000000000000000000";
              \$v2000\ := "00000000000000000000000000000000";
              \$v2001\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 2;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v1999\ & "0001" & \$v2000\ & "0001" & \$v2001\;
              \state\ <= pause_setI2002;
            end if;
          when pause_setII2017 =>
            \$arr1697_ptr_take\(0) := '0';
            \$v2012\ := \$arr1697_ptr_take\;
            if \$v2012\(0) = '1' then
              \state\ <= q_wait2011;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v2006\ := "00000000000000000000000000000000";
              \$v2007\ := "00000000000000000000000000000000";
              \$v2008\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 1;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v2006\ & "0001" & \$v2007\ & "0001" & \$v2008\;
              \state\ <= pause_setI2009;
            end if;
          when pause_setII2021 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2019\ := \$arr1697_ptr_take\;
            if \$v2019\(0) = '1' then
              \state\ <= q_wait2018;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v2013\ := "00000000000000000000000000000000";
              \$v2014\ := "00000000000000000000000000000000";
              \$v2015\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 0;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v2013\ & "0001" & \$v2014\ & "0001" & \$v2015\;
              \state\ <= pause_setI2016;
            end if;
          when pause_setII2025 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2023\ := \$arr1704_ptr_take\;
            if \$v2023\(0) = '1' then
              \state\ <= q_wait2022;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 5;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI2020;
            end if;
          when pause_setII2029 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2027\ := \$arr1704_ptr_take\;
            if \$v2027\(0) = '1' then
              \state\ <= q_wait2026;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 4;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI2024;
            end if;
          when pause_setII2033 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2031\ := \$arr1704_ptr_take\;
            if \$v2031\(0) = '1' then
              \state\ <= q_wait2030;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 3;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI2028;
            end if;
          when pause_setII2037 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2035\ := \$arr1704_ptr_take\;
            if \$v2035\(0) = '1' then
              \state\ <= q_wait2034;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 2;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2032;
            end if;
          when pause_setII2041 =>
            \$arr1704_ptr_take\(0) := '0';
            \$v2039\ := \$arr1704_ptr_take\;
            if \$v2039\(0) = '1' then
              \state\ <= q_wait2038;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 1;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI2036;
            end if;
          when pause_setII2045 =>
            \$arr1703_ptr_take\(0) := '0';
            \$v2043\ := \$arr1704_ptr_take\;
            if \$v2043\(0) = '1' then
              \state\ <= q_wait2042;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 0;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= X"000000" & X"14";
              \state\ <= pause_setI2040;
            end if;
          when pause_setII2049 =>
            \$arr1702_ptr_take\(0) := '0';
            \$v2047\ := \$arr1703_ptr_take\;
            if \$v2047\(0) = '1' then
              \state\ <= q_wait2046;
            else
              \$arr1703_ptr_take\(0) := '1';
              \$arr1703_ptr_write\ <= 0;
              \$arr1703_write_request\ <= '1';
              \$arr1703_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI2044;
            end if;
          when pause_setII2053 =>
            \$arr1701_ptr_take\(0) := '0';
            \$v2051\ := \$arr1702_ptr_take\;
            if \$v2051\(0) = '1' then
              \state\ <= q_wait2050;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2048;
            end if;
          when pause_setII2057 =>
            \$arr1700_ptr_take\(0) := '0';
            \$v2055\ := \$arr1701_ptr_take\;
            if \$v2055\(0) = '1' then
              \state\ <= q_wait2054;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2052;
            end if;
          when pause_setII2061 =>
            \$arr1699_ptr_take\(0) := '0';
            \$v2059\ := \$arr1700_ptr_take\;
            if \$v2059\(0) = '1' then
              \state\ <= q_wait2058;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr_write\ <= 0;
              \$arr1700_write_request\ <= '1';
              \$arr1700_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2056;
            end if;
          when pause_setII2065 =>
            \$arr1698_ptr_take\(0) := '0';
            \$v2063\ := \$arr1699_ptr_take\;
            if \$v2063\(0) = '1' then
              \state\ <= q_wait2062;
            else
              \$arr1699_ptr_take\(0) := '1';
              \$arr1699_ptr_write\ <= 0;
              \$arr1699_write_request\ <= '1';
              \$arr1699_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2060;
            end if;
          when q_wait1714 =>
            \$v1715\ := \$arr1697_ptr_take\;
            if \$v1715\(0) = '1' then
              \state\ <= q_wait1714;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
              \state\ <= pause_getI1712;
            end if;
          when q_wait1718 =>
            \$v1719\ := \$arr1697_ptr_take\;
            if \$v1719\(0) = '1' then
              \state\ <= q_wait1718;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
              \state\ <= pause_getI1716;
            end if;
          when q_wait1726 =>
            \$v1727\ := \$arr1697_ptr_take\;
            if \$v1727\(0) = '1' then
              \state\ <= q_wait1726;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(list_tail700_arg(0 to 31)));
              \state\ <= pause_getI1724;
            end if;
          when q_wait1732 =>
            \$v1733\ := \$arr1702_ptr_take\;
            if \$v1733\(0) = '1' then
              \state\ <= q_wait1732;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= \$325\;
              \state\ <= pause_setI1730;
            end if;
          when q_wait1736 =>
            \$v1737\ := \$arr1702_ptr_take\;
            if \$v1737\(0) = '1' then
              \state\ <= q_wait1736;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1734;
            end if;
          when q_wait1740 =>
            \$v1741\ := \$arr1696_ptr_take\;
            if \$v1741\(0) = '1' then
              \state\ <= q_wait1740;
            else
              \$arr1696_ptr_take\(0) := '1';
              \$arr1696_ptr\ <= to_integer(unsigned(\$328\));
              \state\ <= pause_getI1738;
            end if;
          when q_wait1744 =>
            \$v1745\ := \$arr1702_ptr_take\;
            if \$v1745\(0) = '1' then
              \state\ <= q_wait1744;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1742;
            end if;
          when q_wait1748 =>
            \$v1749\ := \$arr1700_ptr_take\;
            if \$v1749\(0) = '1' then
              \state\ <= q_wait1748;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1746;
            end if;
          when q_wait1752 =>
            \$v1753\ := \$arr1701_ptr_take\;
            if \$v1753\(0) = '1' then
              \state\ <= q_wait1752;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$260_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1750;
            end if;
          when q_wait1759 =>
            \$v1760\ := \$arr1697_ptr_take\;
            if \$v1760\(0) = '1' then
              \state\ <= q_wait1759;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1754\ := eclat_add(\$259_x\ & "00000000000000000000000000000010");
              \$v1755\ := "00000000000000000000000000000000";
              \$v1756\ := "00000000000000000000000000000000";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$260_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1754\ & "0001" & \$v1755\ & "0001" & \$v1756\;
              \state\ <= pause_setI1757;
            end if;
          when q_wait1763 =>
            \$v1764\ := \$arr1701_ptr_take\;
            if \$v1764\(0) = '1' then
              \state\ <= q_wait1763;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$260_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1761;
            end if;
          when q_wait1767 =>
            \$v1768\ := \$arr1697_ptr_take\;
            if \$v1768\(0) = '1' then
              \state\ <= q_wait1767;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$260_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= \$265\;
              \state\ <= pause_setI1765;
            end if;
          when q_wait1773 =>
            \$v1774\ := \$arr1701_ptr_take\;
            if \$v1774\(0) = '1' then
              \state\ <= q_wait1773;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1771;
            end if;
          when q_wait1778 =>
            \$v1779\ := \$arr1701_ptr_take\;
            if \$v1779\(0) = '1' then
              \state\ <= q_wait1778;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1776;
            end if;
          when q_wait1787 =>
            \$v1788\ := \$arr1701_ptr_take\;
            if \$v1788\(0) = '1' then
              \state\ <= q_wait1787;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1785;
            end if;
          when q_wait1791 =>
            \$v1792\ := \$arr1700_ptr_take\;
            if \$v1792\(0) = '1' then
              \state\ <= q_wait1791;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1789;
            end if;
          when q_wait1798 =>
            \$v1799\ := \$arr1697_ptr_take\;
            if \$v1799\(0) = '1' then
              \state\ <= q_wait1798;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1793\ := "00000000000000000000000000000011";
              \$v1794\ := "00000000000000000000000000000000";
              \$v1795\ := "00000000000000000000000000000010";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$279_i\ & "00000000000000000000000000000010")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1793\ & "0001" & \$v1794\ & "0001" & \$v1795\;
              \state\ <= pause_setI1796;
            end if;
          when q_wait1805 =>
            \$v1806\ := \$arr1697_ptr_take\;
            if \$v1806\(0) = '1' then
              \state\ <= q_wait1805;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1800\ := "00000000000000000000000000000011";
              \$v1801\ := eclat_add(\$279_i\ & "00000000000000000000000000000001");
              \$v1802\ := "00000000000000000000000000000010";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$279_i\ & "00000000000000000000000000000010")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1800\ & "0010" & \$v1801\ & "0001" & \$v1802\;
              \state\ <= pause_setI1803;
            end if;
          when q_wait1811 =>
            \$v1812\ := \$arr1701_ptr_take\;
            if \$v1812\(0) = '1' then
              \state\ <= q_wait1811;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1809;
            end if;
          when q_wait1815 =>
            \$v1816\ := \$arr1700_ptr_take\;
            if \$v1816\(0) = '1' then
              \state\ <= q_wait1815;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1813;
            end if;
          when q_wait1820 =>
            \$v1821\ := \$arr1697_ptr_take\;
            if \$v1821\(0) = '1' then
              \state\ <= q_wait1820;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1817\ := "00000000000000000000000000000011";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$288_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & loop3732_arg & "0001" & \$258_len\ & "0001" & \$v1817\;
              \state\ <= pause_setI1818;
            end if;
          when q_wait1825 =>
            \$v1826\ := \$arr1701_ptr_take\;
            if \$v1826\(0) = '1' then
              \state\ <= q_wait1825;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1823;
            end if;
          when q_wait1829 =>
            \$v1830\ := \$arr1700_ptr_take\;
            if \$v1830\(0) = '1' then
              \state\ <= q_wait1829;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1827;
            end if;
          when q_wait1835 =>
            \$v1836\ := \$arr1697_ptr_take\;
            if \$v1836\(0) = '1' then
              \state\ <= q_wait1835;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
              \state\ <= pause_getI1833;
            end if;
          when q_wait1847 =>
            \$v1848\ := \$arr1697_ptr_take\;
            if \$v1848\(0) = '1' then
              \state\ <= q_wait1847;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(loop3732_arg));
              \state\ <= pause_getI1845;
            end if;
          when q_wait1851 =>
            \$v1852\ := \$arr1701_ptr_take\;
            if \$v1852\(0) = '1' then
              \state\ <= q_wait1851;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$84_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1849;
            end if;
          when q_wait1858 =>
            \$v1859\ := \$arr1697_ptr_take\;
            if \$v1859\(0) = '1' then
              \state\ <= q_wait1858;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1853\ := eclat_add(\$76_x\ & "00000000000000000000000000000010");
              \$v1854\ := "00000000000000000000000000000000";
              \$v1855\ := "00000000000000000000000000000000";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$84_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1853\ & "0001" & \$v1854\ & "0001" & \$v1855\;
              \state\ <= pause_setI1856;
            end if;
          when q_wait1862 =>
            \$v1863\ := \$arr1701_ptr_take\;
            if \$v1863\(0) = '1' then
              \state\ <= q_wait1862;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= eclat_add(\$84_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1860;
            end if;
          when q_wait1866 =>
            \$v1867\ := \$arr1697_ptr_take\;
            if \$v1867\(0) = '1' then
              \state\ <= q_wait1866;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$84_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= \$v151\;
              \state\ <= pause_setI1864;
            end if;
          when q_wait1872 =>
            \$v1873\ := \$arr1701_ptr_take\;
            if \$v1873\(0) = '1' then
              \state\ <= q_wait1872;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1870;
            end if;
          when q_wait1877 =>
            \$v1878\ := \$arr1701_ptr_take\;
            if \$v1878\(0) = '1' then
              \state\ <= q_wait1877;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1875;
            end if;
          when q_wait1886 =>
            \$v1887\ := \$arr1701_ptr_take\;
            if \$v1887\(0) = '1' then
              \state\ <= q_wait1886;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1884;
            end if;
          when q_wait1890 =>
            \$v1891\ := \$arr1700_ptr_take\;
            if \$v1891\(0) = '1' then
              \state\ <= q_wait1890;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1888;
            end if;
          when q_wait1897 =>
            \$v1898\ := \$arr1697_ptr_take\;
            if \$v1898\(0) = '1' then
              \state\ <= q_wait1897;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1892\ := "00000000000000000000000000000011";
              \$v1893\ := "00000000000000000000000000000000";
              \$v1894\ := "00000000000000000000000000000010";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$87_i\ & "00000000000000000000000000000010")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1892\ & "0001" & \$v1893\ & "0001" & \$v1894\;
              \state\ <= pause_setI1895;
            end if;
          when q_wait1904 =>
            \$v1905\ := \$arr1697_ptr_take\;
            if \$v1905\(0) = '1' then
              \state\ <= q_wait1904;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1899\ := "00000000000000000000000000000011";
              \$v1900\ := eclat_add(\$87_i\ & "00000000000000000000000000000001");
              \$v1901\ := "00000000000000000000000000000010";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$87_i\ & "00000000000000000000000000000010")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1899\ & "0010" & \$v1900\ & "0001" & \$v1901\;
              \state\ <= pause_setI1902;
            end if;
          when q_wait1910 =>
            \$v1911\ := \$arr1701_ptr_take\;
            if \$v1911\(0) = '1' then
              \state\ <= q_wait1910;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1908;
            end if;
          when q_wait1914 =>
            \$v1915\ := \$arr1700_ptr_take\;
            if \$v1915\(0) = '1' then
              \state\ <= q_wait1914;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1912;
            end if;
          when q_wait1919 =>
            \$v1920\ := \$arr1697_ptr_take\;
            if \$v1920\(0) = '1' then
              \state\ <= q_wait1919;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1916\ := "00000000000000000000000000000011";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$89_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & loop3732_arg & "0001" & len & "0001" & \$v1916\;
              \state\ <= pause_setI1917;
            end if;
          when q_wait1924 =>
            \$v1925\ := \$arr1701_ptr_take\;
            if \$v1925\(0) = '1' then
              \state\ <= q_wait1924;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1922;
            end if;
          when q_wait1928 =>
            \$v1929\ := \$arr1700_ptr_take\;
            if \$v1929\(0) = '1' then
              \state\ <= q_wait1928;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1926;
            end if;
          when q_wait1934 =>
            \$v1935\ := \$arr1697_ptr_take\;
            if \$v1935\(0) = '1' then
              \state\ <= q_wait1934;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(\$220_i\));
              \state\ <= pause_getI1932;
            end if;
          when q_wait1946 =>
            \$v1947\ := \$arr1697_ptr_take\;
            if \$v1947\(0) = '1' then
              \state\ <= q_wait1946;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$arr1697_ptr\ <= to_integer(unsigned(loop3732_arg));
              \state\ <= pause_getI1944;
            end if;
          when q_wait1950 =>
            \$v1951\ := \$arr1700_ptr_take\;
            if \$v1951\(0) = '1' then
              \state\ <= q_wait1950;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1948;
            end if;
          when q_wait1954 =>
            \$v1955\ := \$arr1700_ptr_take\;
            if \$v1955\(0) = '1' then
              \state\ <= q_wait1954;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr_write\ <= 0;
              \$arr1700_write_request\ <= '1';
              \$arr1700_write\ <= eclat_add(\$74_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI1952;
            end if;
          when q_wait1959 =>
            \$v1960\ := \$arr1697_ptr_take\;
            if \$v1960\(0) = '1' then
              \state\ <= q_wait1959;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1956\ := "00000000000000000000000000000000";
              \$arr1697_ptr_write\ <= to_integer(unsigned(eclat_add(\$74_i\ & "00000000000000000000000000000001")));
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$71_x\ & "0010" & loop3732_arg & "0001" & \$v1956\;
              \state\ <= pause_setI1957;
            end if;
          when q_wait1964 =>
            \$v1965\ := \$arr1700_ptr_take\;
            if \$v1965\(0) = '1' then
              \state\ <= q_wait1964;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr\ <= 0;
              \state\ <= pause_getI1962;
            end if;
          when q_wait1968 =>
            \$v1969\ := \$arr1701_ptr_take\;
            if \$v1969\(0) = '1' then
              \state\ <= q_wait1968;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr\ <= 0;
              \state\ <= pause_getI1966;
            end if;
          when q_wait1974 =>
            \$v1975\ := \$arr1702_ptr_take\;
            if \$v1975\(0) = '1' then
              \state\ <= q_wait1974;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= \$v114\;
              \state\ <= pause_setI1972;
            end if;
          when q_wait1978 =>
            \$v1979\ := \$arr1702_ptr_take\;
            if \$v1979\(0) = '1' then
              \state\ <= q_wait1978;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1976;
            end if;
          when q_wait1982 =>
            \$v1983\ := \$arr1696_ptr_take\;
            if \$v1983\(0) = '1' then
              \state\ <= q_wait1982;
            else
              \$arr1696_ptr_take\(0) := '1';
              \$arr1696_ptr\ <= to_integer(unsigned(\$v111\));
              \state\ <= pause_getI1980;
            end if;
          when q_wait1986 =>
            \$v1987\ := \$arr1702_ptr_take\;
            if \$v1987\(0) = '1' then
              \state\ <= q_wait1986;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr\ <= 0;
              \state\ <= pause_getI1984;
            end if;
          when q_wait1990 =>
            \$v1991\ := \$arr1701_ptr_take\;
            if \$v1991\(0) = '1' then
              \state\ <= q_wait1990;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= "00000000000000000000000000000011";
              \state\ <= pause_setI1988;
            end if;
          when q_wait1997 =>
            \$v1998\ := \$arr1697_ptr_take\;
            if \$v1998\(0) = '1' then
              \state\ <= q_wait1997;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1992\ := "00000000000000000000000000000001";
              \$v1993\ := "00000000000000000000000000000010";
              \$v1994\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 3;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0010" & \$v1992\ & "0010" & \$v1993\ & "0001" & \$v1994\;
              \state\ <= pause_setI1995;
            end if;
          when q_wait2004 =>
            \$v2005\ := \$arr1697_ptr_take\;
            if \$v2005\(0) = '1' then
              \state\ <= q_wait2004;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v1999\ := "00000000000000000000000000000000";
              \$v2000\ := "00000000000000000000000000000000";
              \$v2001\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 2;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v1999\ & "0001" & \$v2000\ & "0001" & \$v2001\;
              \state\ <= pause_setI2002;
            end if;
          when q_wait2011 =>
            \$v2012\ := \$arr1697_ptr_take\;
            if \$v2012\(0) = '1' then
              \state\ <= q_wait2011;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v2006\ := "00000000000000000000000000000000";
              \$v2007\ := "00000000000000000000000000000000";
              \$v2008\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 1;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v2006\ & "0001" & \$v2007\ & "0001" & \$v2008\;
              \state\ <= pause_setI2009;
            end if;
          when q_wait2018 =>
            \$v2019\ := \$arr1697_ptr_take\;
            if \$v2019\(0) = '1' then
              \state\ <= q_wait2018;
            else
              \$arr1697_ptr_take\(0) := '1';
              \$v2013\ := "00000000000000000000000000000000";
              \$v2014\ := "00000000000000000000000000000000";
              \$v2015\ := "00000000000000000000000000000101";
              \$arr1697_ptr_write\ <= 0;
              \$arr1697_write_request\ <= '1';
              \$arr1697_write\ <= "0001" & \$v2013\ & "0001" & \$v2014\ & "0001" & \$v2015\;
              \state\ <= pause_setI2016;
            end if;
          when q_wait2022 =>
            \$v2023\ := \$arr1704_ptr_take\;
            if \$v2023\(0) = '1' then
              \state\ <= q_wait2022;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 5;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI2020;
            end if;
          when q_wait2026 =>
            \$v2027\ := \$arr1704_ptr_take\;
            if \$v2027\(0) = '1' then
              \state\ <= q_wait2026;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 4;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI2024;
            end if;
          when q_wait2030 =>
            \$v2031\ := \$arr1704_ptr_take\;
            if \$v2031\(0) = '1' then
              \state\ <= q_wait2030;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 3;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI2028;
            end if;
          when q_wait2034 =>
            \$v2035\ := \$arr1704_ptr_take\;
            if \$v2035\(0) = '1' then
              \state\ <= q_wait2034;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 2;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2032;
            end if;
          when q_wait2038 =>
            \$v2039\ := \$arr1704_ptr_take\;
            if \$v2039\(0) = '1' then
              \state\ <= q_wait2038;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 1;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI2036;
            end if;
          when q_wait2042 =>
            \$v2043\ := \$arr1704_ptr_take\;
            if \$v2043\(0) = '1' then
              \state\ <= q_wait2042;
            else
              \$arr1704_ptr_take\(0) := '1';
              \$arr1704_ptr_write\ <= 0;
              \$arr1704_write_request\ <= '1';
              \$arr1704_write\ <= X"000000" & X"14";
              \state\ <= pause_setI2040;
            end if;
          when q_wait2046 =>
            \$v2047\ := \$arr1703_ptr_take\;
            if \$v2047\(0) = '1' then
              \state\ <= q_wait2046;
            else
              \$arr1703_ptr_take\(0) := '1';
              \$arr1703_ptr_write\ <= 0;
              \$arr1703_write_request\ <= '1';
              \$arr1703_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI2044;
            end if;
          when q_wait2050 =>
            \$v2051\ := \$arr1702_ptr_take\;
            if \$v2051\(0) = '1' then
              \state\ <= q_wait2050;
            else
              \$arr1702_ptr_take\(0) := '1';
              \$arr1702_ptr_write\ <= 0;
              \$arr1702_write_request\ <= '1';
              \$arr1702_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2048;
            end if;
          when q_wait2054 =>
            \$v2055\ := \$arr1701_ptr_take\;
            if \$v2055\(0) = '1' then
              \state\ <= q_wait2054;
            else
              \$arr1701_ptr_take\(0) := '1';
              \$arr1701_ptr_write\ <= 0;
              \$arr1701_write_request\ <= '1';
              \$arr1701_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2052;
            end if;
          when q_wait2058 =>
            \$v2059\ := \$arr1700_ptr_take\;
            if \$v2059\(0) = '1' then
              \state\ <= q_wait2058;
            else
              \$arr1700_ptr_take\(0) := '1';
              \$arr1700_ptr_write\ <= 0;
              \$arr1700_write_request\ <= '1';
              \$arr1700_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2056;
            end if;
          when q_wait2062 =>
            \$v2063\ := \$arr1699_ptr_take\;
            if \$v2063\(0) = '1' then
              \state\ <= q_wait2062;
            else
              \$arr1699_ptr_take\(0) := '1';
              \$arr1699_ptr_write\ <= 0;
              \$arr1699_write_request\ <= '1';
              \$arr1699_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI2060;
            end if;
          when q_wait2066 =>
            \$v2067\ := \$arr1698_ptr_take\;
            if \$v2067\(0) = '1' then
              \state\ <= q_wait2066;
            else
              \$arr1698_ptr_take\(0) := '1';
              \$arr1698_ptr_write\ <= 0;
              \$arr1698_write_request\ <= '1';
              \$arr1698_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI2064;
            end if;
          when compute1707 =>
            rdy1706 := eclat_false;
            \$v2067\ := \$arr1698_ptr_take\;
            if \$v2067\(0) = '1' then
              \state\ <= q_wait2066;
            else
              \$arr1698_ptr_take\(0) := '1';
              \$arr1698_ptr_write\ <= 0;
              \$arr1698_write_request\ <= '1';
              \$arr1698_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI2064;
            end if;
          end case;
          
          result <= result1705;
          rdy <= rdy1706;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
