-- code generated from the following source code:
--   ../RibbitVm/fail.ecl
--   ../RibbitVm/vm.ecl
--
-- with the following command:
--
--    ./eclat ../RibbitVm/fail.ecl ../RibbitVm/vm.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute1456, \$147_forever1811388\, \$147_forever1811389\, \$147_forever1811390\, \$147_forever1811391\, \$147_forever1811392\, \$147_forever1811393\, \$147_forever1811394\, \$147_forever1811395\, \$147_forever1811396\, \$147_forever1811397\, \$147_forever1811398\, \$147_forever1811399\, \$147_forever1811400\, \$147_forever1811401\, \$147_forever1811402\, \$147_forever1811403\, \$147_forever1811404\, \$147_forever1811405\, \$147_forever1811406\, \$147_forever1811407\, \$147_forever1811408\, \$147_forever1811409\, \$147_forever1811410\, \$147_forever1811411\, \$147_forever1811412\, \$147_forever1811413\, \$147_forever1811414\, \$147_forever1811415\, \$147_forever1811416\, \$147_forever1811417\, \$147_forever1811418\, \$147_forever1811419\, \$147_forever1811420\, \$147_forever1811421\, \$147_forever1811422\, \$147_forever1811423\, \$147_forever1811424\, \$147_forever1811425\, \$147_forever1811426\, \$147_forever1811427\, \$147_forever1811428\, \$147_forever1811429\, \$147_forever1811430\, \$147_forever1811431\, \$147_forever1811432\, \$147_forever1811433\, \$147_forever1811434\, \$147_forever1811435\, \$147_forever1811436\, \$147_forever1811437\, \$147_forever1811438\, \$147_forever1811439\, \$147_forever1811440\, \$147_forever1811441\, \$147_forever1811442\, \$147_forever1811443\, \$147_forever1811444\, \$147_forever1811445\, \$147_forever1811446\, \$147_forever1811447\, \$147_forever1811448\, \$147_forever1811449\, \$147_forever1811450\, get_pause1462, get_pause1479, get_pause1504, get_pause1572, get_pause1644, get_pause1661, get_pause1686, get_pause1754, get_pause1826, get_pause1843, get_pause1868, get_pause1936, get_pause2008, get_pause2025, get_pause2050, get_pause2118, get_pause2190, get_pause2206, get_pause2241, get_pause2309, get_pause2381, get_pause2397, get_pause2435, get_pause2503, get_pause2575, get_pause2585, get_pause2615, get_pause2683, get_pause2755, get_pause2765, get_pause2795, get_pause2863, get_pause2935, get_pause2945, get_pause2975, get_pause3043, get_pause3115, get_pause3132, get_pause3157, get_pause3229, get_pause3246, get_pause3271, get_pause3343, get_pause3360, get_pause3385, get_pause3457, get_pause3467, get_pause3499, get_pause3571, get_pause3582, get_pause3622, get_pause3694, get_pause3711, get_pause3729, get_pause3797, get_pause3869, get_pause3886, get_pause3904, get_pause3976, get_pause3986, get_pause4009, get_pause4077, get_pause4145, get_wait1461, get_wait1463, get_wait1478, get_wait1491, get_wait1503, get_wait1512, get_wait1530, get_wait1539, get_wait1544, get_wait1557, get_wait1566, get_wait1571, get_wait1580, get_wait1598, get_wait1607, get_wait1612, get_wait1625, get_wait1634, get_wait1643, get_wait1645, get_wait1660, get_wait1673, get_wait1685, get_wait1694, get_wait1712, get_wait1721, get_wait1726, get_wait1739, get_wait1748, get_wait1753, get_wait1762, get_wait1780, get_wait1789, get_wait1794, get_wait1807, get_wait1816, get_wait1825, get_wait1827, get_wait1842, get_wait1855, get_wait1867, get_wait1876, get_wait1894, get_wait1903, get_wait1908, get_wait1921, get_wait1930, get_wait1935, get_wait1944, get_wait1962, get_wait1971, get_wait1976, get_wait1989, get_wait1998, get_wait2007, get_wait2009, get_wait2024, get_wait2037, get_wait2049, get_wait2058, get_wait2076, get_wait2085, get_wait2090, get_wait2103, get_wait2112, get_wait2117, get_wait2126, get_wait2144, get_wait2153, get_wait2158, get_wait2171, get_wait2180, get_wait2189, get_wait2205, get_wait2229, get_wait2240, get_wait2249, get_wait2267, get_wait2276, get_wait2281, get_wait2294, get_wait2303, get_wait2308, get_wait2317, get_wait2335, get_wait2344, get_wait2349, get_wait2362, get_wait2371, get_wait2380, get_wait2396, get_wait2420, get_wait2434, get_wait2443, get_wait2461, get_wait2470, get_wait2475, get_wait2488, get_wait2497, get_wait2502, get_wait2511, get_wait2529, get_wait2538, get_wait2543, get_wait2556, get_wait2565, get_wait2574, get_wait2584, get_wait2602, get_wait2614, get_wait2623, get_wait2641, get_wait2650, get_wait2655, get_wait2668, get_wait2677, get_wait2682, get_wait2691, get_wait2709, get_wait2718, get_wait2723, get_wait2736, get_wait2745, get_wait2754, get_wait2764, get_wait2782, get_wait2794, get_wait2803, get_wait2821, get_wait2830, get_wait2835, get_wait2848, get_wait2857, get_wait2862, get_wait2871, get_wait2889, get_wait2898, get_wait2903, get_wait2916, get_wait2925, get_wait2934, get_wait2944, get_wait2962, get_wait2974, get_wait2983, get_wait3001, get_wait3010, get_wait3015, get_wait3028, get_wait3037, get_wait3042, get_wait3051, get_wait3069, get_wait3078, get_wait3083, get_wait3096, get_wait3105, get_wait3114, get_wait3116, get_wait3131, get_wait3144, get_wait3156, get_wait3165, get_wait3183, get_wait3192, get_wait3197, get_wait3210, get_wait3219, get_wait3228, get_wait3230, get_wait3245, get_wait3258, get_wait3270, get_wait3279, get_wait3297, get_wait3306, get_wait3311, get_wait3324, get_wait3333, get_wait3342, get_wait3344, get_wait3359, get_wait3372, get_wait3384, get_wait3393, get_wait3411, get_wait3420, get_wait3425, get_wait3438, get_wait3447, get_wait3456, get_wait3466, get_wait3484, get_wait3498, get_wait3507, get_wait3525, get_wait3534, get_wait3539, get_wait3552, get_wait3561, get_wait3570, get_wait3581, get_wait3600, get_wait3609, get_wait3621, get_wait3630, get_wait3648, get_wait3657, get_wait3662, get_wait3675, get_wait3684, get_wait3693, get_wait3695, get_wait3710, get_wait3723, get_wait3728, get_wait3737, get_wait3755, get_wait3764, get_wait3769, get_wait3782, get_wait3791, get_wait3796, get_wait3805, get_wait3823, get_wait3832, get_wait3837, get_wait3850, get_wait3859, get_wait3868, get_wait3870, get_wait3885, get_wait3898, get_wait3903, get_wait3912, get_wait3930, get_wait3939, get_wait3944, get_wait3957, get_wait3966, get_wait3975, get_wait3985, get_wait4003, get_wait4008, get_wait4017, get_wait4035, get_wait4044, get_wait4049, get_wait4062, get_wait4071, get_wait4076, get_wait4085, get_wait4103, get_wait4112, get_wait4117, get_wait4130, get_wait4139, get_wait4144, get_wait4153, get_wait4171, get_wait4180, get_wait4185, get_wait4198, get_wait4207, get_wait4216, pause_getI1464, pause_getI1468, pause_getI1480, pause_getI1492, pause_getI1508, pause_getI1513, pause_getI1517, pause_getI1526, pause_getI1531, pause_getI1535, pause_getI1540, pause_getI1545, pause_getI1553, pause_getI1558, pause_getI1562, pause_getI1567, pause_getI1576, pause_getI1581, pause_getI1585, pause_getI1594, pause_getI1599, pause_getI1603, pause_getI1608, pause_getI1613, pause_getI1621, pause_getI1626, pause_getI1630, pause_getI1635, pause_getI1646, pause_getI1650, pause_getI1662, pause_getI1674, pause_getI1690, pause_getI1695, pause_getI1699, pause_getI1708, pause_getI1713, pause_getI1717, pause_getI1722, pause_getI1727, pause_getI1735, pause_getI1740, pause_getI1744, pause_getI1749, pause_getI1758, pause_getI1763, pause_getI1767, pause_getI1776, pause_getI1781, pause_getI1785, pause_getI1790, pause_getI1795, pause_getI1803, pause_getI1808, pause_getI1812, pause_getI1817, pause_getI1828, pause_getI1832, pause_getI1844, pause_getI1856, pause_getI1872, pause_getI1877, pause_getI1881, pause_getI1890, pause_getI1895, pause_getI1899, pause_getI1904, pause_getI1909, pause_getI1917, pause_getI1922, pause_getI1926, pause_getI1931, pause_getI1940, pause_getI1945, pause_getI1949, pause_getI1958, pause_getI1963, pause_getI1967, pause_getI1972, pause_getI1977, pause_getI1985, pause_getI1990, pause_getI1994, pause_getI1999, pause_getI2010, pause_getI2014, pause_getI2026, pause_getI2038, pause_getI2054, pause_getI2059, pause_getI2063, pause_getI2072, pause_getI2077, pause_getI2081, pause_getI2086, pause_getI2091, pause_getI2099, pause_getI2104, pause_getI2108, pause_getI2113, pause_getI2122, pause_getI2127, pause_getI2131, pause_getI2140, pause_getI2145, pause_getI2149, pause_getI2154, pause_getI2159, pause_getI2167, pause_getI2172, pause_getI2176, pause_getI2181, pause_getI2191, pause_getI2207, pause_getI2230, pause_getI2245, pause_getI2250, pause_getI2254, pause_getI2263, pause_getI2268, pause_getI2272, pause_getI2277, pause_getI2282, pause_getI2290, pause_getI2295, pause_getI2299, pause_getI2304, pause_getI2313, pause_getI2318, pause_getI2322, pause_getI2331, pause_getI2336, pause_getI2340, pause_getI2345, pause_getI2350, pause_getI2358, pause_getI2363, pause_getI2367, pause_getI2372, pause_getI2382, pause_getI2398, pause_getI2421, pause_getI2439, pause_getI2444, pause_getI2448, pause_getI2457, pause_getI2462, pause_getI2466, pause_getI2471, pause_getI2476, pause_getI2484, pause_getI2489, pause_getI2493, pause_getI2498, pause_getI2507, pause_getI2512, pause_getI2516, pause_getI2525, pause_getI2530, pause_getI2534, pause_getI2539, pause_getI2544, pause_getI2552, pause_getI2557, pause_getI2561, pause_getI2566, pause_getI2576, pause_getI2586, pause_getI2603, pause_getI2608, pause_getI2619, pause_getI2624, pause_getI2628, pause_getI2637, pause_getI2642, pause_getI2646, pause_getI2651, pause_getI2656, pause_getI2664, pause_getI2669, pause_getI2673, pause_getI2678, pause_getI2687, pause_getI2692, pause_getI2696, pause_getI2705, pause_getI2710, pause_getI2714, pause_getI2719, pause_getI2724, pause_getI2732, pause_getI2737, pause_getI2741, pause_getI2746, pause_getI2756, pause_getI2766, pause_getI2783, pause_getI2788, pause_getI2799, pause_getI2804, pause_getI2808, pause_getI2817, pause_getI2822, pause_getI2826, pause_getI2831, pause_getI2836, pause_getI2844, pause_getI2849, pause_getI2853, pause_getI2858, pause_getI2867, pause_getI2872, pause_getI2876, pause_getI2885, pause_getI2890, pause_getI2894, pause_getI2899, pause_getI2904, pause_getI2912, pause_getI2917, pause_getI2921, pause_getI2926, pause_getI2936, pause_getI2946, pause_getI2963, pause_getI2968, pause_getI2979, pause_getI2984, pause_getI2988, pause_getI2997, pause_getI3002, pause_getI3006, pause_getI3011, pause_getI3016, pause_getI3024, pause_getI3029, pause_getI3033, pause_getI3038, pause_getI3047, pause_getI3052, pause_getI3056, pause_getI3065, pause_getI3070, pause_getI3074, pause_getI3079, pause_getI3084, pause_getI3092, pause_getI3097, pause_getI3101, pause_getI3106, pause_getI3117, pause_getI3121, pause_getI3133, pause_getI3145, pause_getI3150, pause_getI3161, pause_getI3166, pause_getI3170, pause_getI3179, pause_getI3184, pause_getI3188, pause_getI3193, pause_getI3198, pause_getI3206, pause_getI3211, pause_getI3215, pause_getI3220, pause_getI3231, pause_getI3235, pause_getI3247, pause_getI3259, pause_getI3264, pause_getI3275, pause_getI3280, pause_getI3284, pause_getI3293, pause_getI3298, pause_getI3302, pause_getI3307, pause_getI3312, pause_getI3320, pause_getI3325, pause_getI3329, pause_getI3334, pause_getI3345, pause_getI3349, pause_getI3361, pause_getI3373, pause_getI3378, pause_getI3389, pause_getI3394, pause_getI3398, pause_getI3407, pause_getI3412, pause_getI3416, pause_getI3421, pause_getI3426, pause_getI3434, pause_getI3439, pause_getI3443, pause_getI3448, pause_getI3458, pause_getI3468, pause_getI3485, pause_getI3503, pause_getI3508, pause_getI3512, pause_getI3521, pause_getI3526, pause_getI3530, pause_getI3535, pause_getI3540, pause_getI3548, pause_getI3553, pause_getI3557, pause_getI3562, pause_getI3572, pause_getI3583, pause_getI3601, pause_getI3605, pause_getI3610, pause_getI3615, pause_getI3626, pause_getI3631, pause_getI3635, pause_getI3644, pause_getI3649, pause_getI3653, pause_getI3658, pause_getI3663, pause_getI3671, pause_getI3676, pause_getI3680, pause_getI3685, pause_getI3696, pause_getI3700, pause_getI3712, pause_getI3724, pause_getI3733, pause_getI3738, pause_getI3742, pause_getI3751, pause_getI3756, pause_getI3760, pause_getI3765, pause_getI3770, pause_getI3778, pause_getI3783, pause_getI3787, pause_getI3792, pause_getI3801, pause_getI3806, pause_getI3810, pause_getI3819, pause_getI3824, pause_getI3828, pause_getI3833, pause_getI3838, pause_getI3846, pause_getI3851, pause_getI3855, pause_getI3860, pause_getI3871, pause_getI3875, pause_getI3887, pause_getI3899, pause_getI3908, pause_getI3913, pause_getI3917, pause_getI3926, pause_getI3931, pause_getI3935, pause_getI3940, pause_getI3945, pause_getI3953, pause_getI3958, pause_getI3962, pause_getI3967, pause_getI3977, pause_getI3987, pause_getI4004, pause_getI4013, pause_getI4018, pause_getI4022, pause_getI4031, pause_getI4036, pause_getI4040, pause_getI4045, pause_getI4050, pause_getI4058, pause_getI4063, pause_getI4067, pause_getI4072, pause_getI4081, pause_getI4086, pause_getI4090, pause_getI4099, pause_getI4104, pause_getI4108, pause_getI4113, pause_getI4118, pause_getI4126, pause_getI4131, pause_getI4135, pause_getI4140, pause_getI4149, pause_getI4154, pause_getI4158, pause_getI4167, pause_getI4172, pause_getI4176, pause_getI4181, pause_getI4186, pause_getI4194, pause_getI4199, pause_getI4203, pause_getI4208, pause_getI4212, pause_getI4217, pause_getII1465, pause_getII1469, pause_getII1481, pause_getII1493, pause_getII1509, pause_getII1514, pause_getII1518, pause_getII1527, pause_getII1532, pause_getII1536, pause_getII1541, pause_getII1546, pause_getII1554, pause_getII1559, pause_getII1563, pause_getII1568, pause_getII1577, pause_getII1582, pause_getII1586, pause_getII1595, pause_getII1600, pause_getII1604, pause_getII1609, pause_getII1614, pause_getII1622, pause_getII1627, pause_getII1631, pause_getII1636, pause_getII1647, pause_getII1651, pause_getII1663, pause_getII1675, pause_getII1691, pause_getII1696, pause_getII1700, pause_getII1709, pause_getII1714, pause_getII1718, pause_getII1723, pause_getII1728, pause_getII1736, pause_getII1741, pause_getII1745, pause_getII1750, pause_getII1759, pause_getII1764, pause_getII1768, pause_getII1777, pause_getII1782, pause_getII1786, pause_getII1791, pause_getII1796, pause_getII1804, pause_getII1809, pause_getII1813, pause_getII1818, pause_getII1829, pause_getII1833, pause_getII1845, pause_getII1857, pause_getII1873, pause_getII1878, pause_getII1882, pause_getII1891, pause_getII1896, pause_getII1900, pause_getII1905, pause_getII1910, pause_getII1918, pause_getII1923, pause_getII1927, pause_getII1932, pause_getII1941, pause_getII1946, pause_getII1950, pause_getII1959, pause_getII1964, pause_getII1968, pause_getII1973, pause_getII1978, pause_getII1986, pause_getII1991, pause_getII1995, pause_getII2000, pause_getII2011, pause_getII2015, pause_getII2027, pause_getII2039, pause_getII2055, pause_getII2060, pause_getII2064, pause_getII2073, pause_getII2078, pause_getII2082, pause_getII2087, pause_getII2092, pause_getII2100, pause_getII2105, pause_getII2109, pause_getII2114, pause_getII2123, pause_getII2128, pause_getII2132, pause_getII2141, pause_getII2146, pause_getII2150, pause_getII2155, pause_getII2160, pause_getII2168, pause_getII2173, pause_getII2177, pause_getII2182, pause_getII2192, pause_getII2208, pause_getII2231, pause_getII2246, pause_getII2251, pause_getII2255, pause_getII2264, pause_getII2269, pause_getII2273, pause_getII2278, pause_getII2283, pause_getII2291, pause_getII2296, pause_getII2300, pause_getII2305, pause_getII2314, pause_getII2319, pause_getII2323, pause_getII2332, pause_getII2337, pause_getII2341, pause_getII2346, pause_getII2351, pause_getII2359, pause_getII2364, pause_getII2368, pause_getII2373, pause_getII2383, pause_getII2399, pause_getII2422, pause_getII2440, pause_getII2445, pause_getII2449, pause_getII2458, pause_getII2463, pause_getII2467, pause_getII2472, pause_getII2477, pause_getII2485, pause_getII2490, pause_getII2494, pause_getII2499, pause_getII2508, pause_getII2513, pause_getII2517, pause_getII2526, pause_getII2531, pause_getII2535, pause_getII2540, pause_getII2545, pause_getII2553, pause_getII2558, pause_getII2562, pause_getII2567, pause_getII2577, pause_getII2587, pause_getII2604, pause_getII2609, pause_getII2620, pause_getII2625, pause_getII2629, pause_getII2638, pause_getII2643, pause_getII2647, pause_getII2652, pause_getII2657, pause_getII2665, pause_getII2670, pause_getII2674, pause_getII2679, pause_getII2688, pause_getII2693, pause_getII2697, pause_getII2706, pause_getII2711, pause_getII2715, pause_getII2720, pause_getII2725, pause_getII2733, pause_getII2738, pause_getII2742, pause_getII2747, pause_getII2757, pause_getII2767, pause_getII2784, pause_getII2789, pause_getII2800, pause_getII2805, pause_getII2809, pause_getII2818, pause_getII2823, pause_getII2827, pause_getII2832, pause_getII2837, pause_getII2845, pause_getII2850, pause_getII2854, pause_getII2859, pause_getII2868, pause_getII2873, pause_getII2877, pause_getII2886, pause_getII2891, pause_getII2895, pause_getII2900, pause_getII2905, pause_getII2913, pause_getII2918, pause_getII2922, pause_getII2927, pause_getII2937, pause_getII2947, pause_getII2964, pause_getII2969, pause_getII2980, pause_getII2985, pause_getII2989, pause_getII2998, pause_getII3003, pause_getII3007, pause_getII3012, pause_getII3017, pause_getII3025, pause_getII3030, pause_getII3034, pause_getII3039, pause_getII3048, pause_getII3053, pause_getII3057, pause_getII3066, pause_getII3071, pause_getII3075, pause_getII3080, pause_getII3085, pause_getII3093, pause_getII3098, pause_getII3102, pause_getII3107, pause_getII3118, pause_getII3122, pause_getII3134, pause_getII3146, pause_getII3151, pause_getII3162, pause_getII3167, pause_getII3171, pause_getII3180, pause_getII3185, pause_getII3189, pause_getII3194, pause_getII3199, pause_getII3207, pause_getII3212, pause_getII3216, pause_getII3221, pause_getII3232, pause_getII3236, pause_getII3248, pause_getII3260, pause_getII3265, pause_getII3276, pause_getII3281, pause_getII3285, pause_getII3294, pause_getII3299, pause_getII3303, pause_getII3308, pause_getII3313, pause_getII3321, pause_getII3326, pause_getII3330, pause_getII3335, pause_getII3346, pause_getII3350, pause_getII3362, pause_getII3374, pause_getII3379, pause_getII3390, pause_getII3395, pause_getII3399, pause_getII3408, pause_getII3413, pause_getII3417, pause_getII3422, pause_getII3427, pause_getII3435, pause_getII3440, pause_getII3444, pause_getII3449, pause_getII3459, pause_getII3469, pause_getII3486, pause_getII3504, pause_getII3509, pause_getII3513, pause_getII3522, pause_getII3527, pause_getII3531, pause_getII3536, pause_getII3541, pause_getII3549, pause_getII3554, pause_getII3558, pause_getII3563, pause_getII3573, pause_getII3584, pause_getII3602, pause_getII3606, pause_getII3611, pause_getII3616, pause_getII3627, pause_getII3632, pause_getII3636, pause_getII3645, pause_getII3650, pause_getII3654, pause_getII3659, pause_getII3664, pause_getII3672, pause_getII3677, pause_getII3681, pause_getII3686, pause_getII3697, pause_getII3701, pause_getII3713, pause_getII3725, pause_getII3734, pause_getII3739, pause_getII3743, pause_getII3752, pause_getII3757, pause_getII3761, pause_getII3766, pause_getII3771, pause_getII3779, pause_getII3784, pause_getII3788, pause_getII3793, pause_getII3802, pause_getII3807, pause_getII3811, pause_getII3820, pause_getII3825, pause_getII3829, pause_getII3834, pause_getII3839, pause_getII3847, pause_getII3852, pause_getII3856, pause_getII3861, pause_getII3872, pause_getII3876, pause_getII3888, pause_getII3900, pause_getII3909, pause_getII3914, pause_getII3918, pause_getII3927, pause_getII3932, pause_getII3936, pause_getII3941, pause_getII3946, pause_getII3954, pause_getII3959, pause_getII3963, pause_getII3968, pause_getII3978, pause_getII3988, pause_getII4005, pause_getII4014, pause_getII4019, pause_getII4023, pause_getII4032, pause_getII4037, pause_getII4041, pause_getII4046, pause_getII4051, pause_getII4059, pause_getII4064, pause_getII4068, pause_getII4073, pause_getII4082, pause_getII4087, pause_getII4091, pause_getII4100, pause_getII4105, pause_getII4109, pause_getII4114, pause_getII4119, pause_getII4127, pause_getII4132, pause_getII4136, pause_getII4141, pause_getII4150, pause_getII4155, pause_getII4159, pause_getII4168, pause_getII4173, pause_getII4177, pause_getII4182, pause_getII4187, pause_getII4195, pause_getII4200, pause_getII4204, pause_getII4209, pause_getII4213, pause_getII4218, pause_setI1457, pause_setI1474, pause_setI1485, pause_setI1521, pause_setI1589, pause_setI1639, pause_setI1656, pause_setI1667, pause_setI1703, pause_setI1771, pause_setI1821, pause_setI1838, pause_setI1849, pause_setI1885, pause_setI1953, pause_setI2003, pause_setI2020, pause_setI2031, pause_setI2067, pause_setI2135, pause_setI2185, pause_setI2201, pause_setI2213, pause_setI2223, pause_setI2258, pause_setI2326, pause_setI2376, pause_setI2392, pause_setI2404, pause_setI2414, pause_setI2452, pause_setI2520, pause_setI2570, pause_setI2580, pause_setI2592, pause_setI2596, pause_setI2632, pause_setI2700, pause_setI2750, pause_setI2760, pause_setI2772, pause_setI2776, pause_setI2812, pause_setI2880, pause_setI2930, pause_setI2940, pause_setI2952, pause_setI2956, pause_setI2992, pause_setI3060, pause_setI3110, pause_setI3127, pause_setI3138, pause_setI3174, pause_setI3224, pause_setI3241, pause_setI3252, pause_setI3288, pause_setI3338, pause_setI3355, pause_setI3366, pause_setI3402, pause_setI3452, pause_setI3462, pause_setI3474, pause_setI3478, pause_setI3516, pause_setI3566, pause_setI3577, pause_setI3589, pause_setI3594, pause_setI3639, pause_setI3689, pause_setI3706, pause_setI3717, pause_setI3746, pause_setI3814, pause_setI3864, pause_setI3881, pause_setI3892, pause_setI3921, pause_setI3971, pause_setI3981, pause_setI3993, pause_setI3997, pause_setI4026, pause_setI4094, pause_setI4162, pause_setI4221, pause_setI4225, pause_setI4229, pause_setI4233, pause_setI4237, pause_setII1458, pause_setII1475, pause_setII1486, pause_setII1522, pause_setII1590, pause_setII1640, pause_setII1657, pause_setII1668, pause_setII1704, pause_setII1772, pause_setII1822, pause_setII1839, pause_setII1850, pause_setII1886, pause_setII1954, pause_setII2004, pause_setII2021, pause_setII2032, pause_setII2068, pause_setII2136, pause_setII2186, pause_setII2202, pause_setII2214, pause_setII2224, pause_setII2259, pause_setII2327, pause_setII2377, pause_setII2393, pause_setII2405, pause_setII2415, pause_setII2453, pause_setII2521, pause_setII2571, pause_setII2581, pause_setII2593, pause_setII2597, pause_setII2633, pause_setII2701, pause_setII2751, pause_setII2761, pause_setII2773, pause_setII2777, pause_setII2813, pause_setII2881, pause_setII2931, pause_setII2941, pause_setII2953, pause_setII2957, pause_setII2993, pause_setII3061, pause_setII3111, pause_setII3128, pause_setII3139, pause_setII3175, pause_setII3225, pause_setII3242, pause_setII3253, pause_setII3289, pause_setII3339, pause_setII3356, pause_setII3367, pause_setII3403, pause_setII3453, pause_setII3463, pause_setII3475, pause_setII3479, pause_setII3517, pause_setII3567, pause_setII3578, pause_setII3590, pause_setII3595, pause_setII3640, pause_setII3690, pause_setII3707, pause_setII3718, pause_setII3747, pause_setII3815, pause_setII3865, pause_setII3882, pause_setII3893, pause_setII3922, pause_setII3972, pause_setII3982, pause_setII3994, pause_setII3998, pause_setII4027, pause_setII4095, pause_setII4163, pause_setII4222, pause_setII4226, pause_setII4230, pause_setII4234, pause_setII4238, q_wait1459, q_wait1466, q_wait1470, q_wait1476, q_wait1482, q_wait1487, q_wait1494, q_wait1510, q_wait1515, q_wait1519, q_wait1523, q_wait1528, q_wait1533, q_wait1537, q_wait1542, q_wait1547, q_wait1555, q_wait1560, q_wait1564, q_wait1569, q_wait1578, q_wait1583, q_wait1587, q_wait1591, q_wait1596, q_wait1601, q_wait1605, q_wait1610, q_wait1615, q_wait1623, q_wait1628, q_wait1632, q_wait1637, q_wait1641, q_wait1648, q_wait1652, q_wait1658, q_wait1664, q_wait1669, q_wait1676, q_wait1692, q_wait1697, q_wait1701, q_wait1705, q_wait1710, q_wait1715, q_wait1719, q_wait1724, q_wait1729, q_wait1737, q_wait1742, q_wait1746, q_wait1751, q_wait1760, q_wait1765, q_wait1769, q_wait1773, q_wait1778, q_wait1783, q_wait1787, q_wait1792, q_wait1797, q_wait1805, q_wait1810, q_wait1814, q_wait1819, q_wait1823, q_wait1830, q_wait1834, q_wait1840, q_wait1846, q_wait1851, q_wait1858, q_wait1874, q_wait1879, q_wait1883, q_wait1887, q_wait1892, q_wait1897, q_wait1901, q_wait1906, q_wait1911, q_wait1919, q_wait1924, q_wait1928, q_wait1933, q_wait1942, q_wait1947, q_wait1951, q_wait1955, q_wait1960, q_wait1965, q_wait1969, q_wait1974, q_wait1979, q_wait1987, q_wait1992, q_wait1996, q_wait2001, q_wait2005, q_wait2012, q_wait2016, q_wait2022, q_wait2028, q_wait2033, q_wait2040, q_wait2056, q_wait2061, q_wait2065, q_wait2069, q_wait2074, q_wait2079, q_wait2083, q_wait2088, q_wait2093, q_wait2101, q_wait2106, q_wait2110, q_wait2115, q_wait2124, q_wait2129, q_wait2133, q_wait2137, q_wait2142, q_wait2147, q_wait2151, q_wait2156, q_wait2161, q_wait2169, q_wait2174, q_wait2178, q_wait2183, q_wait2187, q_wait2193, q_wait2203, q_wait2209, q_wait2215, q_wait2225, q_wait2232, q_wait2247, q_wait2252, q_wait2256, q_wait2260, q_wait2265, q_wait2270, q_wait2274, q_wait2279, q_wait2284, q_wait2292, q_wait2297, q_wait2301, q_wait2306, q_wait2315, q_wait2320, q_wait2324, q_wait2328, q_wait2333, q_wait2338, q_wait2342, q_wait2347, q_wait2352, q_wait2360, q_wait2365, q_wait2369, q_wait2374, q_wait2378, q_wait2384, q_wait2394, q_wait2400, q_wait2406, q_wait2416, q_wait2423, q_wait2441, q_wait2446, q_wait2450, q_wait2454, q_wait2459, q_wait2464, q_wait2468, q_wait2473, q_wait2478, q_wait2486, q_wait2491, q_wait2495, q_wait2500, q_wait2509, q_wait2514, q_wait2518, q_wait2522, q_wait2527, q_wait2532, q_wait2536, q_wait2541, q_wait2546, q_wait2554, q_wait2559, q_wait2563, q_wait2568, q_wait2572, q_wait2578, q_wait2582, q_wait2588, q_wait2594, q_wait2598, q_wait2605, q_wait2610, q_wait2621, q_wait2626, q_wait2630, q_wait2634, q_wait2639, q_wait2644, q_wait2648, q_wait2653, q_wait2658, q_wait2666, q_wait2671, q_wait2675, q_wait2680, q_wait2689, q_wait2694, q_wait2698, q_wait2702, q_wait2707, q_wait2712, q_wait2716, q_wait2721, q_wait2726, q_wait2734, q_wait2739, q_wait2743, q_wait2748, q_wait2752, q_wait2758, q_wait2762, q_wait2768, q_wait2774, q_wait2778, q_wait2785, q_wait2790, q_wait2801, q_wait2806, q_wait2810, q_wait2814, q_wait2819, q_wait2824, q_wait2828, q_wait2833, q_wait2838, q_wait2846, q_wait2851, q_wait2855, q_wait2860, q_wait2869, q_wait2874, q_wait2878, q_wait2882, q_wait2887, q_wait2892, q_wait2896, q_wait2901, q_wait2906, q_wait2914, q_wait2919, q_wait2923, q_wait2928, q_wait2932, q_wait2938, q_wait2942, q_wait2948, q_wait2954, q_wait2958, q_wait2965, q_wait2970, q_wait2981, q_wait2986, q_wait2990, q_wait2994, q_wait2999, q_wait3004, q_wait3008, q_wait3013, q_wait3018, q_wait3026, q_wait3031, q_wait3035, q_wait3040, q_wait3049, q_wait3054, q_wait3058, q_wait3062, q_wait3067, q_wait3072, q_wait3076, q_wait3081, q_wait3086, q_wait3094, q_wait3099, q_wait3103, q_wait3108, q_wait3112, q_wait3119, q_wait3123, q_wait3129, q_wait3135, q_wait3140, q_wait3147, q_wait3152, q_wait3163, q_wait3168, q_wait3172, q_wait3176, q_wait3181, q_wait3186, q_wait3190, q_wait3195, q_wait3200, q_wait3208, q_wait3213, q_wait3217, q_wait3222, q_wait3226, q_wait3233, q_wait3237, q_wait3243, q_wait3249, q_wait3254, q_wait3261, q_wait3266, q_wait3277, q_wait3282, q_wait3286, q_wait3290, q_wait3295, q_wait3300, q_wait3304, q_wait3309, q_wait3314, q_wait3322, q_wait3327, q_wait3331, q_wait3336, q_wait3340, q_wait3347, q_wait3351, q_wait3357, q_wait3363, q_wait3368, q_wait3375, q_wait3380, q_wait3391, q_wait3396, q_wait3400, q_wait3404, q_wait3409, q_wait3414, q_wait3418, q_wait3423, q_wait3428, q_wait3436, q_wait3441, q_wait3445, q_wait3450, q_wait3454, q_wait3460, q_wait3464, q_wait3470, q_wait3476, q_wait3480, q_wait3487, q_wait3505, q_wait3510, q_wait3514, q_wait3518, q_wait3523, q_wait3528, q_wait3532, q_wait3537, q_wait3542, q_wait3550, q_wait3555, q_wait3559, q_wait3564, q_wait3568, q_wait3574, q_wait3579, q_wait3585, q_wait3591, q_wait3596, q_wait3603, q_wait3607, q_wait3612, q_wait3617, q_wait3628, q_wait3633, q_wait3637, q_wait3641, q_wait3646, q_wait3651, q_wait3655, q_wait3660, q_wait3665, q_wait3673, q_wait3678, q_wait3682, q_wait3687, q_wait3691, q_wait3698, q_wait3702, q_wait3708, q_wait3714, q_wait3719, q_wait3726, q_wait3735, q_wait3740, q_wait3744, q_wait3748, q_wait3753, q_wait3758, q_wait3762, q_wait3767, q_wait3772, q_wait3780, q_wait3785, q_wait3789, q_wait3794, q_wait3803, q_wait3808, q_wait3812, q_wait3816, q_wait3821, q_wait3826, q_wait3830, q_wait3835, q_wait3840, q_wait3848, q_wait3853, q_wait3857, q_wait3862, q_wait3866, q_wait3873, q_wait3877, q_wait3883, q_wait3889, q_wait3894, q_wait3901, q_wait3910, q_wait3915, q_wait3919, q_wait3923, q_wait3928, q_wait3933, q_wait3937, q_wait3942, q_wait3947, q_wait3955, q_wait3960, q_wait3964, q_wait3969, q_wait3973, q_wait3979, q_wait3983, q_wait3989, q_wait3995, q_wait3999, q_wait4006, q_wait4015, q_wait4020, q_wait4024, q_wait4028, q_wait4033, q_wait4038, q_wait4042, q_wait4047, q_wait4052, q_wait4060, q_wait4065, q_wait4069, q_wait4074, q_wait4083, q_wait4088, q_wait4092, q_wait4096, q_wait4101, q_wait4106, q_wait4110, q_wait4115, q_wait4120, q_wait4128, q_wait4133, q_wait4137, q_wait4142, q_wait4151, q_wait4156, q_wait4160, q_wait4164, q_wait4169, q_wait4174, q_wait4178, q_wait4183, q_wait4188, q_wait4196, q_wait4201, q_wait4205, q_wait4210, q_wait4214, q_wait4219, q_wait4223, q_wait4227, q_wait4231, q_wait4235, q_wait4239);
  signal \state\: t_state;
  type array_value_1 is array (natural range <>) of value(0 to 0);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  type array_value_108 is array (natural range <>) of value(0 to 107);
  signal arr1451 : array_value_108(0 to 89999) := (others => (others => '0'));
  signal \$arr1451_value\ : value(0 to 107);
  signal \$arr1451_ptr\ : natural range 0 to 89999;
  signal \$arr1451_ptr_write\ : natural range 0 to 89999;
  signal \$arr1451_write\ : value(0 to 107);
  signal \$arr1451_write_request\ : std_logic := '0';
  signal arr1452 : array_value_32(0 to 4) := (others => (others => '0'));
  signal \$arr1452_value\ : value(0 to 31);
  signal \$arr1452_ptr\ : natural range 0 to 4;
  signal \$arr1452_ptr_write\ : natural range 0 to 4;
  signal \$arr1452_write\ : value(0 to 31);
  signal \$arr1452_write_request\ : std_logic := '0';
  signal arr1453 : array_value_1(0 to 19) := (others => (others => '0'));
  signal \$arr1453_value\ : value(0 to 0);
  signal \$arr1453_ptr\ : natural range 0 to 19;
  signal \$arr1453_ptr_write\ : natural range 0 to 19;
  signal \$arr1453_write\ : value(0 to 0);
  signal \$arr1453_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1451_write_request\ = '1' then
                    arr1451(\$arr1451_ptr_write\) <= \$arr1451_write\;
                  else
                   \$arr1451_value\ <= arr1451(\$arr1451_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1452_write_request\ = '1' then
                    arr1452(\$arr1452_ptr_write\) <= \$arr1452_write\;
                  else
                   \$arr1452_value\ <= arr1452(\$arr1452_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1453_write_request\ = '1' then
                    arr1453(\$arr1453_ptr_write\) <= \$arr1453_write\;
                  else
                   \$arr1453_value\ <= arr1453(\$arr1453_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$814\, \$v3432\, \$v2617\, \$v2482\, \$v1938\, \$1396_x\, 
               \$411\, \$v2730\, \$1153\, \$825\, \$1302\, \$193\, \$v2097\, 
               \$v2052\, \$v1574\, \$v1863\, \$70_y\, \$1463\, \$1573\, 
               \$1520\, \$839_x\, \$v2910\, \$v1915\, \$752\, \$v1551\, 
               \$888\, \$354\, \$446\, \$709\, \$v4056\, \$860\, \$v1681\, 
               \$v2977\, \$1274\, \$166\, \$426_y\, \$1111\, \$v2236\, 
               \$1552_x\, \$1342\, \$270_x\, \$1630\, \$v1870\, \$v3268\, 
               \$v1501\, \$v3731\, \$365\, \$v1801\, \$v3204\, \$v2243\, 
               \$969\, \$590\, \$337\, \$1270_x\, \$425_x\, \$1341\, 
               \$v4124\, \$1556\, \$797\, \$997\, \$v2437\, \$v2972\, 
               \$632_x\, \$1504\, \$688_x\, \$692\, \$224_x\, \$v2612\, 
               \$v3022\, \$1016\, \$v3624\, \$877\, \$316_x\, \$948_x\, 
               \$1100\, \$633_y\, \$1665\, \$274\, \$v3090\, \$1291\, \$291\, 
               \$540_x\, \$v2047\, \$338\, \$318_result_after_f\, \$v3273\, 
               \$1083\, \$463\, \$492\, \$165\, \$333_x\, \$83_x\, \$v25\, 
               \$v2238\, \$v3318\, \$v3844\, \$646\, \$986\, \$902_x\, 
               \$1152\, \$v2797\, \$v2311\, \$209_result_after_f\, \$v4192\, 
               \$245\, \$1446\, \$1332_x\, \$379_x\, \$1648\, \$442_x\, 
               \$71_result_after_f\, \$663\, \$1602\, \$1079_x\, \$793_x\, 
               \$v3045\, \$v3496\, \$768\, \$1531\, \$561\, \$v2288\, 
               \$1221\, \$447\, \$1603\, \$v2550\, \$1358\, \$934\, \$642_x\, 
               \$v2505\, \$1238\, \$400\, \$1275\, \$674\, \$76_result\, 
               \$161_x\, \$275\, \$v2120\, \$v3951\, \$65_x\, \$906\, \$798\, 
               \$1212_x\, \$73_result\, \$v35\, \$720\, \$v3546\, \$55_x\, 
               \$v3501\, \$208_y\, \$520\, \$851_x\, \$1143_x\, \$53_y\, 
               \$v4147\, \$1337_x\, \$1222\, \$207_x\, \$v3619\, \$v3776\, 
               \$1011_x\, \$1249\, \$1428\, \$v3159\, \$1598_x\, \$1148_x\, 
               \$v3387\, \$v2685\, \$v2045\, \$1401\, \$1169\, \$693\, 
               \$1400\, \$1032\, \$v2662\, \$v1688\, \$v1683\, \$302\, 
               \$v3799\, \$v4011\, \$1584\, \$586_x\, \$v2792\, \$317_y\, 
               \$1676\, \$v3906\, \$1503\, \$256\, \$1369\, \$v1865\, \$923\, 
               \$v2427\, \$779\, \$1447\, \$v2842\, \$1217_x\, \$v1506\, 
               \$427_result_after_f\, \$1043\, \$182\, \$67_z\, \$488_x\, 
               \$545\, \$v42\, \$v1619\, \$1383_x\, \$v2165\, \$1644_x\, 
               \$1442_x\, \$965_x\, \$84_x\, \$v2356\, \$66_y\, \$1619\, 
               \$v2430\, \$1499_x\, \$509\, \$383\, \$1474\, \$960_x\, 
               \$970\, \$1649\, \$52_x\, \$v3154\, \$607\, \$61_y\, \$856_x\, 
               \$1557\, \$591\, \$747_x\, \$v1733\, \$618\, \$493\, \$v2432\, 
               \$69_x\, \$572\, \$v3382\, \$474\, \$v36\, \$647\, \$v3669\, 
               \$544\, \$1015\, \$1074_x\, \$v1756\, \$751\, \$1180\, 
               \$v1499\, \$228\, \$v2865\, \$v1983\, \$384\, \$907\, 
               \$v4079\, \$229\, \$1084\, \$1417\, \$861\ : value(0 to 35) := (others => '0');
      variable \$1067\, \$1136\, \$1392\, \$1495\, \$v75\, \$326\, \$1205\, 
               \$435\, \$217\ : value(0 to 63) := (others => '0');
      variable \$v1916\, \$v2731\, \$v3502\, \$v1871\, \$v2312\, \$v1757\, 
               \$v2686\, \$v4080\, \$v4012\, \$v3155\, \$v3952\, \$v3620\, 
               \$v2438\, \$v3845\, \$v3497\, \$v3274\, \$v2237\, \$v2433\, 
               \$v3269\, \$v1682\, \$v2121\, \$v1500\, \$v3160\, \$v3732\, 
               \$v2973\, \$v2046\, \$v2551\, \$v1866\, \$v1507\, \$v4057\, 
               \$v2911\, \$v2166\, \$v2239\, \$v2048\, \$v2244\, \$v1689\, 
               \$v2289\, \$v1734\, \$v1620\, \$v1939\, \$v3205\, \$v2053\, 
               \$v3670\, \$v2098\, \$v2978\, \$v3625\, \$v2843\, \$v3777\, 
               \$v2663\, \$v2793\, \$v3383\, \$v3023\, \$v3907\, \$v2431\, 
               \$v1984\, \$v3319\, \$v1802\, \$v2866\, \$v2798\, \$v3046\, 
               \$v2483\, \$v4148\, \$v1684\, \$v1575\, \$v3091\, \$v1864\, 
               \$v3547\, \$v4125\, \$v2506\, \$v4193\, \$v2428\, \$v3800\, 
               \$v2613\, \$v2618\, \$v1552\, \$v1502\, \$v3433\, \$v2357\, 
               \$v3388\ : value(0 to 3) := (others => '0');
      variable \$v2501\, \$v98\, \$867_lock\, \$v39_lock\, \$v1698\, 
               \$v1556\, \$v2379\, \$v1611\, \$887_lock\, \$1166_lock\, 
               \$192_lock\, \$1538_lock\, \$v3019\, \$1010_lock\, \$v2075\, 
               \$v2210\, \$v2660\, \$v3287\, \$v1672\, \$1130_lock\, 
               \$453_lock\, \$1236_lock\, \$v2474\, \$v97\, \$179_lock\, 
               \$846_lock\, \$v3849\, \$1235_lock\, \$v3674\, \$804_lock\, 
               \$v2095\, \$1281_lock\, \$v3055\, \$v2080\, \$v4152\, 
               \$v1592\, \$v2227\, \$v2339\, \$661_lock\, \$533_lock\, 
               \$1315_lock\, \$505_lock\, \$215_lock\, \$764_lock\, \$v3878\, 
               \$v2879\, \$v2542\, \$1159_lock\, \$v3332\, \$v1975\, 
               \$v4228\, \$242_lock\, \$1427_lock\, \$v2649\, \$1262_lock\, 
               \$v3934\, \$v1602\, \$v1543\, \$v2699\, \$499_lock\, 
               \$778_lock\, \$v3173\, \$v3519\, \$v2573\, \$v2920\, \$v102\, 
               \$v2834\, \$1218\, \$v4007\, \$v2961\, \$v4220\, \$v1725\, 
               \$v1716\, \$v3727\, \$489\, \$v3143\, \$v1934\, \$v1617\, 
               \$v3817\, \$v58_lock\, \$v2325\, \$v4138\, \$v2908\, \$v3397\, 
               \$v1835\, \$v2157\, \$v4175\, \$v2515\, \$1616_lock\, 
               \$v1925\, \$v4070\, \$v1970\, \$1510_lock\, \$v1888\, 
               \$v1665\, \$v1649\, \$v1477\, \$v4093\, \$v1766\, \$983_lock\, 
               \$v2194\, \$v4039\, \$1617_lock\, \$v2759\, \$v2966\, 
               \$481_lock\, \$1683_lock\, \$v1907\, \$1583_lock\, 
               \$1118_lock\, \$v2455\, \$v2667\, \$v4061\, \$v2717\, 
               \$v2070\, \$v1495\, \$921_lock\, \$v2595\, \$v2460\, \$v3929\, 
               \$919_lock\, \$v1831\, \$v3073\, \$v2407\, \$1615_lock\, 
               \$v2184\, \$v3371\, \$v43_lock\, \$1098_lock\, \$v4157\, 
               \$706_lock\, \$507_lock\, \$1134_lock\, \$v1948\, \$v3560\, 
               \$1394_lock\, \$v3858\, \$344_lock\, \$v1460\, \$351_lock\, 
               \$v2888\, \$v3895\, \$v2321\, \$895_lock\, \$v2672\, 
               \$461_lock\, \$1287_lock\, \$v4001\, \$v1913\, \$901_lock\, 
               \$v3759\, \$378_lock\, \$v2753\, \$v1730\, \$v3938\, \$v2839\, 
               \$v2293\, \$269_lock\, \$v1738\, \$v94\, \$v3911\, \$v3586\, 
               \$v2233\, \$v3608\, \$v3647\, \$315_lock\, \$v3419\, \$v2253\, 
               \$811_lock\, \$v1538\, \$v2695\, \$v1898\, \$v2062\, \$v2479\, 
               \$v2907\, \$v1853\, \$1271\, \$v2955\, \$v2057\, \$v4002\, 
               \$v3316\, \$v1966\, \$v1902\, \$334\, \$v3948\, \$1355_lock\, 
               \$v1774\, \$v60_lock\, \$v3683\, \$v3328\, \$v1824\, \$v2779\, 
               \$v2138\, \$v3656\, \$857\, \$v3341\, \$v3709\, \$v2519\, 
               \$v3182\, \$v1670\, \$v117\, \$v3763\, \$1376_lock\, 
               \$288_lock\, \$v3401\, \$263_lock\, \$v2547\, \$1461_lock\, 
               \$v2640\, \$v4215\, \$v2883\, \$v3688\, \$v2713\, \$v1847\, 
               \$410_lock\, \$v3529\, \$v4232\, \$634_result\, \$v3455\, 
               \$v3446\, \$v1490\, \$v3348\, \$v2353\, \$v3863\, \$v55_lock\, 
               \$845_lock\, \$v2029\, \$v2442\, \$1643_lock\, \$v3703\, 
               \$v2006\, \$v3569\, \$v3148\, \$v22_lock\, \$v2469\, 
               \$1028_lock\, \$v2875\, \$206_lock\, \$1459_lock\, 
               \$1167_lock\, \$v3575\, \$1497_lock\, \$v3679\, \$v1779\, 
               \$639_lock\, \$v3786\, \$v3202\, \$v2564\, \$v3477\, 
               \$605_lock\, \$v1980\, \$v3471\, \$v1884\, \$v3813\, \$v26\, 
               \$v3050\, \$812_lock\, \$v3177\, \$v4066\, \$v2933\, \$v3262\, 
               \$850_lock\, \$432_lock\, \$v3749\, \$1655_lock\, 
               \$1029_lock\, \$1599\, \$v28_lock\, \$1301_lock\, \$v2188\, 
               \$v4075\, \$1570_lock\, \$v3315\, \$v1693\, \$1368_lock\, 
               \$v1929\, \$v4134\, \$v3209\, \$v2375\, \$v3100\, \$v3890\, 
               \$v3027\, \$v4240\, \$459_lock\, \$1637_lock\, \$v4043\, 
               \$v108\, \$v2548\, \$271\, \$1228_lock\, \$v1638\, \$v2861\, 
               \$v1579\, \$1597_lock\, \$v2424\, \$v2763\, \$v2447\, 
               \$v3481\, \$1662_lock\, \$933_lock\, \$941_lock\, \$v31_lock\, 
               \$v2316\, \$v2216\, \$473_lock\, \$v4161\, \$1441_lock\, 
               \$v2162\, \$920_lock\, \$v3009\, \$v3556\, \$1288_lock\, 
               \$235_lock\, \$v2510\, \$v2847\, \$v2987\, \$551_lock\, 
               \$982_lock\, \$v2807\, \$v2924\, \$v2645\, \$v1642\, 
               \$758_lock\, \$1193_lock\, \$v3201\, \$v1720\, \$v2708\, 
               \$v3924\, \$v2606\, \$v1920\, \$v4021\, \$1481_lock\, 
               \$v4016\, \$v3088\, \$v2395\, \$v3358\, \$1493_lock\, 
               \$v2257\, \$v2102\, \$v2840\, \$v4129\, \$200_lock\, \$v2094\, 
               \$v2163\, \$541\, \$v3515\, \$v2960\, \$v3533\, \$v3136\, 
               \$1211_lock\, \$v2939\, \$v2023\, \$v2982\, \$v78_lock\, 
               \$v2528\, \$v4000\, \$287_lock\, \$v3580\, \$v3032\, 
               \$172_lock\, \$v2555\, \$v89\, \$v1584\, \$1397\, \$v4179\, 
               \$v1952\, \$v3506\, \$v114\, \$v2041\, \$v1549\, \$v96\, 
               \$v3305\, \$v1752\, \$v2148\, \$v3142\, \$v4102\, \$v4189\, 
               \$v3692\, \$v3323\, \$1544_lock\, \$v3077\, \$v2690\, 
               \$v2893\, \$913_lock\, \$v3041\, \$v45_lock\, \$v2811\, 
               \$824_lock\, \$955_lock\, \$v73_lock\, \$v1788\, \$v2959\, 
               \$v3482\, \$v2084\, \$v2111\, \$v76_lock\, \$v3278\, \$v1671\, 
               \$380\, \$1661_lock\, \$1187_lock\, \$v4048\, \$v3781\, 
               \$v2722\, \$v4025\, \$v2361\, \$v1561\, \$559_lock\, \$1012\, 
               \$v1981\, \$v2995\, \$v3598\, \$527_lock\, \$v3255\, 
               \$1030_lock\, \$v3005\, \$v2496\, \$1591_lock\, \$v2343\, 
               \$v67_lock\, \$v1880\, \$699_lock\, \$v3296\, \$v3874\, 
               \$v4107\, \$v3667\, \$1530_lock\, \$v104\, \$v2583\, \$v3036\, 
               \$v3538\, \$v2134\, \$v2385\, \$1110_lock\, \$v1943\, result, 
               \$1663_lock\, \$v2035\, \$1645\, \$v1659\, \$v2487\, 
               \$1487_lock\, \$v3842\, \$v1806\, \$v2271\, \$180_lock\, 
               \$1407_lock\, \$v2775\, \$v3613\, \$v1961\, \$v2769\, 
               \$v2820\, \$v1489\, \$v3721\, \$v3773\, \$v2791\, \$v3715\, 
               \$v1633\, \$v3424\, \$v1784\, \$241_lock\, \$v3736\, 
               \$1517_lock\, \$v2781\, \$437_lock\, \$v2066\, \$v2334\, 
               \$v2261\, \$1065_lock\, \$1061_lock\, \$v3376\, \$219_lock\, 
               \$v3916\, \$v3352\, \$v1875\, \$719_lock\, \$v2017\, 
               \$328_lock\, \$v2897\, \$v3381\, \$1269_lock\, \$653_lock\, 
               \$585_lock\, \$v3896\, \$v3227\, \$1550_lock\, \$v1997\, 
               \$v2417\, \$1689_lock\, \$v3902\, \$v3544\, \$v1706\, 
               \$v3661\, \$v2870\, \$v1616\, \$v2635\, \$v1467\, \$v3642\, 
               \$1498_lock\, \$v2589\, \$v3524\, \$1563_lock\, \$1354_lock\, 
               \$1549_lock\, \$v3565\, \$v2579\, \$v1988\, \$1199_lock\, 
               \$1309_lock\, \$418_lock\, \$v3511\, \$631_lock\, \$v2451\, 
               \$748\, \$1338\, \$v1471\, \$v3218\, \$v3283\, \$398_lock\, 
               \$v4202\, \$1096_lock\, \$903\, \$v2002\, \$v2740\, \$966\, 
               \$1453_lock\, \$v3841\, \$487_lock\, \$v3000\, \$1042_lock\, 
               \$v4089\, \$1414_lock\, \$v3191\, \$557_lock\, \$460_lock\, 
               \$875_lock\, \$v2727\, \$v3634\, \$390_lock\, \$v1711\, 
               \$v2601\, \$v2130\, \$v3410\, \$1256_lock\, \$v1677\, 
               \$v2622\, \$v3970\, \$v3465\, \$v3666\, \$996_lock\, \$v1548\, 
               \$1073_lock\, \$v27_lock\, \$v3169\, \$v2815\, \$v2856\, 
               \$324_lock\, \$v3087\, \$v2152\, \$v3543\, \$1165_lock\, 
               \$681_lock\, \$v2659\, \$v3214\, \$v2537\, \$v3291\, \$v1761\, 
               \$v4143\, \$v2654\, \$v3618\, \$v4122\, \$v2929\, \$v2703\, 
               \$v3990\, \$v1852\, \$810_lock\, \$v3961\, \$v1770\, \$v4165\, 
               \$v1811\, \$v4224\, \$243_lock\, \$765_lock\, \$v2802\, 
               \$1629_lock\, \$v3164\, \$323_lock\, \$1149\, \$v3020\, 
               \$v3854\, \$v2465\, \$v3430\, \$v2492\, \$1320_lock\, 
               \$1050_lock\, \$v2902\, \$v2852\, \$v120\, \$v3974\, 
               \$1460_lock\, \$v3301\, \$v2307\, \$v1912\, \$v3187\, 
               \$1609_lock\, \$1389_lock\, \$v3980\, \$v2560\, \$v1653\, 
               \$v1841\, \$587\, \$v2611\, \$v2401\, \$v2116\, \$v3014\, 
               \$v3943\, \$v3082\, \$1473_lock\, \$v2034\, \$1056_lock\, 
               \$v2275\, \$1142_lock\, \$v3442\, \$v3059\, \$v3996\, \$1553\, 
               \$738_lock\, \$v4190\, \$660_lock\, \$v3774\, \$424_lock\, 
               \$1413_lock\, \$v1483\, \$v1993\, \$v3754\, \$v4184\, 
               \$733_lock\, \$v3364\, \$v2266\, \$v2786\, \$v1516\, 
               \$792_lock\, result1454, \$640_lock\, \$v1893\, \$625_lock\, 
               \$v2170\, \$225\, \$372_lock\, \$v1793\, \$1435_lock\, 
               \$v3551\, \$1022_lock\, \$v2735\, \$1518_lock\, rdy1455, 
               \$v3836\, \$v2533\, \$v1629\, \$v2569\, \$v3451\, \$727_lock\, 
               \$976_lock\, \$1004_lock\, \$v2298\, \$v3130\, \$433_lock\, 
               \$v2285\, \$v3223\, \$794\, \$v1743\, \$v4170\, \$v1488\, 
               \$766_lock\, \$v3867\, \$v3405\, \$v91\, \$443\, \$v111\, 
               \$v2370\, \$1289_lock\, \$438_lock\, \$1090_lock\, \$v2107\, 
               \$396_lock\, \$v2627\, \$v3599\, \$603_lock\, \$397_lock\, 
               \$v1520\, \$1179_lock\, \$214_lock\, \$162\, \$v1731\, 
               \$1207_lock\, \$1097_lock\, \$v3238\, \$v1798\, \$558_lock\, 
               \$v2366\, \$v2780\, \$v2523\, \$281_lock\, \$1415_lock\, 
               \$v3415\, \$786_lock\, \$v2728\, \$v4197\, \$v2971\, \$v1747\, 
               \$v3109\, \$v3920\, \$659_lock\, \$v1511\, \$1382_lock\, 
               \$v2013\, \$v3592\, \$641_lock\, \$v3196\, \$832_lock\, 
               \$v2175\, \$v3741\, \$v3153\, \$v3720\, \$579_lock\, \$v4111\, 
               \$v1799\, \$v4236\, \$1234_lock\, \$1324_lock\, \$v2143\, 
               \$1516_lock\, \$v3827\, \$v4097\, \$519_lock\, \$v2480\, 
               \$v4053\, \$v3768\, \$v1854\, \$1551_lock\, \$v3809\, 
               \$v3483\, \$v3629\, \$v3244\, \$v2991\, \$v2248\, \$301_lock\, 
               \$v4121\, \$v2089\, \$v3604\, \$309_lock\, \$v2676\, 
               \$1569_lock\, \$v3429\, \$v1859\, \$v95\, \$v93\, \$604_lock\, 
               \$v3790\, \$v2681\, \$329_lock\, \$v1606\, \$v3392\, \$643\, 
               \$v1524\, \$959_lock\, \$v3884\, \$v3063\, \$1395_lock\, 
               \$1571_lock\, \$v3897\, \$v4116\, \$v106\, \$v2204\, \$v2280\, 
               \$v2036\, \$v3256\, \$352_lock\, \$v2418\, \$838_lock\, 
               \$v3965\, \$873_lock\, \$v2600\, \$v2228\, \$v3831\, \$v3699\, 
               \$v3488\, \$v19_lock\, \$1356_lock\, \$v3250\, \$v3257\, 
               \$v1588\, \$v4054\, \$v2419\, \$1267_lock\, \$v3461\, 
               \$v3822\, \$v3267\, \$v2943\, \$v2329\, \$v4034\, \$v3638\, 
               \$673_lock\, \$v4029\, \$1124_lock\, \$255_lock\, 
               \$1069_lock\, \$743_lock\, \$1268_lock\, \$1443\, \$v2915\, 
               \$707_lock\, \$1675_lock\, \$v3984\, \$v3337\, \$1348_lock\, 
               \$v3068\, \$v2749\, \$617_lock\, \$220_lock\, \$v3597\, 
               \$364_lock\, \$v3437\, \$954_lock\, \$v4084\, \$178_lock\, 
               \$v1529\, \$1248_lock\, \$v2631\, \$v3095\, \$v1956\, 
               \$v2179\, \$1328_lock\, \$1138_lock\, \$v1624\, \$v1820\, 
               \$v1570\, \$v3745\, \$v2354\, \$v3956\, \$v3310\, \$289_lock\, 
               \$v2829\, \$947_lock\, \$v100\, \$v3949\, \$1492_lock\, 
               \$506_lock\, \$687_lock\, \$v3804\, \$v2599\, \$v3369\, 
               \$v2226\, \$v3104\, \$984_lock\, \$v2744\, \$v3234\, \$v2825\, 
               \$v4206\, \$v3120\, \$v3370\, \$1203_lock\, \$v3141\, \$1080\, 
               \$1500\, \$v2348\, \$1390_lock\, \$v1702\, \$v3113\, 
               \$705_lock\, \$v3652\, \$571_lock\, \$v1815\, \$v1597\, 
               \$874_lock\, \$v1534\, \$689\, \$597_lock\, \$v2302\, 
               \$v2125\, \$v4211\, \$v2286\, \$739_lock\, \$v16_lock\, 
               \$v2949\, \$v3124\, \$v3795\, \$v1565\, \$350_lock\, \$v3722\ : value(0 to 0) := (others => '0');
      variable \$1371\, \$1160\, \$345\, \$v18\, \$1684\, \$359\, \$1564\, 
               \$1632\, \$1296\, \$626\, \$819\, \$859\, \$805\, \$589\, 
               \$v24\, \$58_result\, \$1604\, \$1422\, \$v80\, \$773\, 
               \$296\, \$v41\, \$753\, \$1430\, \$1402\, \$339\, \$454\, 
               \$250\, \$528\, \$1343\, \$1154\, \$391\, \$862\, \$799\, 
               \$833\, \$1151\, \$491\, \$1223\, \$1610\, \$1182\, \$1251\, 
               \$1014\, \$552\, \$1188\, \$468\, \$230\, \$612\, \$977\, 
               \$971\, \$195\, \$1276\, \$580\, \$v21\, \$v33\, \$167\, 
               \$1533\, \$908\, \$942\, \$1023\, \$276\, \$905\, \$654\, 
               \$1273\, \$1505\, \$914\, \$694\, \$682\, \$187\, \$1282\, 
               \$1656\, \$1476\, \$1539\, \$882\, \$1082\, \$1511\, \$1113\, 
               \$1377\, \$413\, \$949_y\, \$273\, \$1085\, \$236\, \$1502\, 
               \$1017\, \$310\, \$592\, \$787\, \$574\, \$781\, \$896\, 
               \$1650\, \$676\, \$1454\, \$514\, \$1091\, \$304\, \$367\, 
               \$264\, \$1436\, \$1349\, \$522\, \$373\, \$1647\, \$282\, 
               \$336\, \$796\, \$728\, \$1310\, \$840_y\, \$722\, \$1051\, 
               \$1624\, \$936\, \$448\, \$1005\, \$1340\, \$620\, \$991\, 
               \$405\, \$1037\, \$648\, \$385\, \$645\, \$1555\, \$691\, 
               \$1592\, \$1678\, \$1194_result\, \$1638\, \$173\, \$1578\, 
               \$258\, \$201\, \$1525\, \$1229\, \$1105\, \$999\, \$1586\, 
               \$1363\, \$543\, \$227\, \$1304\, \$1670\, \$1601\, \$928\, 
               \$868\, \$74_result_after_f\, \$v38\, \$714\, \$59_tos\, 
               \$419\, \$56_y\, \$476\, \$668\, \$1045\, \$968\, \$700\, 
               \$1257\, \$1482\, \$598\, \$566\, \$1445\, \$1125_result\, 
               \$1448\, \$164\, \$546\, \$1399\, \$445\, \$1408\, \$482\, 
               \$1174\, \$827\, \$1468\, \$1243\, \$382\, \$v30\, \$750\, 
               \$494\, \$1558\, \$500\, \$1119\, \$759\, \$1220\, \$890\ : value(0 to 107) := (others => '0');
      variable \$1353\, \$1615\, \$v1836\, \$617\, \$1620_i\, \$1355\, 
               \$804\, \$1347\, \$1413\, \$344\, \$178\, \$1544\, \$286\, 
               \$1509\, \$1135\, \$1412\, \$v2607\, \$v2222\, \$680\, 
               \$1394\, \$1543\, \$508\, \$625\, \$1391\, \$329\, \$219\, 
               \$v2524\, \$641\, \$240\, \$1395\, \$1480\, \$635_i\, \$763\, 
               \$409\, \$1124\, \$v3473\, \$570\, \$1280\, \$919\, \$183_i\, 
               \$1487\, \$1496\, \$292_i\, \$1027\, \$734_i\, \$1288\, 
               \$809\, \$v2235\, \$887\, \$1494\, \$v77\, \$1328\, \$1538\, 
               \$v3263\, \$v60\, \$v29\, \$410\, st, \$v3353\, \$v3545\, 
               \$v2310\, \$1666_i\, \$913\, \$v3292\, \$1118\, \$1385_i\, 
               \$v3880\, \$v2389\, \$v4191\, \$396\, \$792\, \$v3879\, 
               \$v2591\, \$901\, \$v1775\, \$395\, \$1435\, \$v1937\, 
               \$v2071\, \$660\, \$459\, \$220\, \$510_i\, \$v2976\, \$262\, 
               \$1600\, \$v2221\, \$813\, \$v3203\, \$v3905\, \$1636\, 
               \$815_i\, \$v2770\, \$878_i\, \$v3089\, \$1021\, \$244\, 
               \$v1496\, \$1309\, \$v1679\, \$v2951\, \$726\, \$791\, \$218\, 
               \$v3623\, \$v3668\, \$767\, \$1654\, \$309\, \$v3818\, 
               \$v2386\, \$v2616\, \$363\, \$1481\, \$v3704\, \$235\, 
               \$v2196\, \$487\, \$v2590\, \$519\, \$v3406\, \$v2864\, 
               \$v1680\, \$1472\, \$630\, \$1572\, \$872\, \$v3775\, 
               \$1574_i\, \$1515\, \$v1666\, \$1123\, \$518\, \$v78\, 
               \$1109\, \$v3044\, \$733\, \$29_a\, \$288\, \$1004\, \$1674\, 
               \$216\, \$246_i\, \$v3158\, \$1583\, \$v1848\, \$1164\, 
               \$900\, \$v3643\, \$1101_i\, \$v2387\, \$v2030\, b, \$397\, 
               \$1434\, \$662\, \$698\, \$1159\, \$1219\, \$v2481\, \$v2436\, 
               \$v2456\, \$1068\, \$1591\, \$1440\, \$v1755\, \$987_i\, 
               \$894\, \$v27\, \$v3489\, \$v3925\, \$922\, \$1590\, \$v1550\, 
               \$v2355\, \$498\, \$967\, \$1545_i\, \$1646\, \$1292_i\, 
               \$831\, \$837\, \$v2412\, \$v19\, \$1227\, \$1643\, \$1234\, 
               \$v2217\, \$417\, \$v3491\, \$v1837\, \$1398\, \$596\, 
               \$1486\, \$1041\, \$280\, \$1186\, \$832\, \$996\, \$371\, 
               \$874\, \$26_a\, \$1211\, \$v2164\, \$v79\, \$841_i\, 
               \$v2199\, \$585\, \$1348\, \$v3239\, \$1090\, \$1089\, 
               \$v2220\, \$v2197\, \$263\, \$578\, \$866\, \$v1862\, \$946\, 
               \$940\, \$1416\, \$1256\, \$137_i\, \$1049\, \$867\, \$v44\, 
               \$924_i\, \$v3493\, \$1057_i\, \$506\, \$v4078\, \$v45\, 
               \$v2051\, \$381\, \$v2841\, \$976\, \$v4010\, \$557\, stbl, 
               \$718\, \$v23\, \$873\, \$179\, \$1126_i\, \$1376\, \$192\, 
               \$v2661\, \$1233\, \$886\, \$424\, ia, \$1427\, \$1682\, 
               \$932\, \$82_i\, \$390\, \$1614\, \$241\, \$v3588\, \$1498\, 
               \$351\, \$v3716\, \$838\, \$v2195\, \$226\, \$v2816\, \$1009\, 
               \$975\, \$v2242\, \$v1593\, \$1314\, \$v3576\, \$1563\, 
               \$1660\, \$1110\, \$1582\, \$v2402\, \$343\, \$769_i\, \$558\, 
               \$v2212\, \$325\, \$1537\, \$1464_i\, \$959\, \$v2429\, 
               \$378\, \$1488_i\, \$353\, \$v3377\, \$v2287\, \$315\, \$v39\, 
               \$1642\, \$v2409\, \$1235\, \$v1861\, \$v2391\, \$v1498\, 
               \$749\, \$858\, \$v2884\, \$743\, \$490\, \$v2411\, \$v4098\, 
               \$551\, \$v2413\, \$1661\, \$1521_i\, \$v2390\, \$v2200\, 
               \$1381\, \$335\, \$v3240\, \$550\, \$603\, \$1597\, \$328\, 
               \$1099\, \$1453\, \$v3843\, \$604\, \$1554\, \$v1655\, \$765\, 
               \$1239_i\, pc, \$v2909\, \$533\, \$631\, \$1683\, \$785\, 
               \$1204\, \$v3520\, \$823\, \$v3587\, \$1367\, \$1066\, 
               \$1042\, \$v17\, \$v2139\, \$777\, \$542\, \$v1525\, \$v3021\, 
               \$1570\, \$v40\, ta, \$v2218\, \$1460\, \$1272\, \$355_i\, 
               \$1142\, \$1003\, \$v3178\, \$1418_i\, \$1688\, \$624\, 
               \$1050\, \$579\, \$608_i\, \$686\, \$v4030\, \$672\, \$527\, 
               \$961_i\, \$1675\, \$1081\, \$1414\, \$v2729\, pos, \$1165\, 
               \$1170_i\, \$652\, \$v1573\, \$673\, \$v2950\, \$1029\, 
               \$v4166\, \$377\, \$995\, \$v4123\, \$1568\, \$v1914\, 
               \$v1860\, \$350\, \$v1732\, \$803\, \$171\, \$1510\, \$1013\, 
               \$1459\, \$269\, \$1301\, \$191\, \$v3365\, \$32_a\, \$v1707\, 
               \$1150\, \$242\, \$1033_i\, \$1179\, \$v73\, \$v1654\, 
               \$v2967\, \$v2234\, \$1444\, \$v3494\, \$423\, \$1664\, 
               \$v16\, \$1290\, \$597\, \$1028\, \$983\, \$458\, \$681\, 
               \$1517\, \$v1678\, \$758\, \$v2410\, \$438\, \$v3492\, \$462\, 
               \$1117\, \$35_a\, \$659\, \$v3593\, \$1359_i\, \$1247\, 
               \$526\, \$933\, \$210_i\, \$1187\, \$1056\, \$1382\, \$255\, 
               \$1096\, \$172\, \$985\, \$v2219\, \$v3490\, \$v3137\, \$481\, 
               \$v1687\, \$135_i\, \$499\, \$v1957\, \$764\, \$319_i\, 
               \$1689\, \$1333_i\, \$v3317\, \$1261\, \$824\, \$v2044\, 
               \$v2425\, \$v3992\, \$1158\, \$v2119\, \$v3730\, \$1458\, 
               \$v1869\, \$199\, \$v2018\, \$1519\, \$v2787\, \$453\, 
               \$v1505\, \$v3500\, \$719\, \$v28\, \$1308\, \$460\, \$300\, 
               \$v1497\, \$181\, \$v3750\, \$v3251\, \$v3472\, \$1315\, 
               \$v3354\, \$616\, \$947\, \$1516\, \$1596\, \$v1800\, 
               \$v2403\, \$v3125\, \$664_i\, \$v1889\, \$v2043\, \$1075_i\, 
               \$1637\, \$1069\, \$v20\, \$428_i\, \$1206\, \$308\, \$1452\, 
               \$1213_i\, \$918\, \$876\, \$v4055\, \$1406\, \$287\, \$920\, 
               \$644\, \$904\, \$504\, \$1662\, \$1616\, \$895\, \$708\, 
               \$1166\, \$v74\, \$1248\, \$v31\, \$v3991\, \$811\, \$1473\, 
               \$v3064\, \$1569\, \$532\, \$1551\, \$706\, \$434\, \$301\, 
               \$1501\, \$505\, \$1609\, \$v2704\, \$399\, \$912\, \$v2796\, 
               \$1137\, \$290\, \$v2426\, \$v3950\, \$v2636\, \$1300\, 
               \$1207\, \$372\, \$1441\, \$1144_i\, \$1192\, \$1629\, \$690\, 
               \$1316_i\, \$786\, \$v2684\, tb, \$v37\, \$1138\, \$1393\, 
               \$602\, \$710_i\, \$584\, \$1368\, \$389\, \$206\, \$1426\, 
               \$v3126\, \$1497\, \$562_i\, \$810\, \$1281\, \$349\, \$437\, 
               \$571\, \$727\, \$687\, \$757\, \$v2096\, \$v4146\, \$852_i\, 
               \$1237\, \$v2042\, \$588\, \$1530\, \$v3614\, \$606\, 
               \$v2211\, \$268\, \$480\, \$v2504\, \$v1618\, \$1269\, \$281\, 
               \$1097\, \$950_i\, \$1655\, \$v1472\, \$v2408\, \$1262\, 
               \$1095\, \$v22\, \$1022\, \$254\, \$1375\, \$732\, \$v2771\, 
               \$560\, \$177\, \$v3149\, \$941\, \$1168\, \$200\, \$778\, 
               \$704\, \$v2262\, \$556\, \$v2330\, \$v3798\, \$1073\, \$982\, 
               \$v2198\, \$81_i\, \$850\, \$1462\, \$v2996\, \$705\, \$v32\, 
               \$1055\, \$795\, \$v1484\, \$314\, \$1010\, \$1031\, \$1608\, 
               \$327\, \$486\, \$1357\, ib, \$364\, \$1286\, \$1255\, 
               \$v2388\, \$163\, \$1193\, \$1263_i\, \$1339\, \$1407\, 
               \$464_i\, \$1287\, \$1354\, \$v3431\, \$v3495\, \$v1473\, 
               \$981\, sp, \$401_i\, \$472\, \$v3705\, \$1618\, \$1529\, 
               \$205\, \$v3386\, \$653\, \$418\, \$v2019\, \$1178\, \$1628\, 
               \$444\, \$452\, \$v3891\, \$1562\, \$436\, \$658\, \$v3272\, 
               \$1195_i\, \$272\, \$v1982\, \$v2549\, \$1228\, a, \$234\, 
               \$473\, \$699\ : value(0 to 31) := (others => '0');
      variable \$arr1451_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1452_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1453_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v3722\); default_zero(\$699\); 
          default_zero(\$350_lock\); default_zero(\$473\); 
          default_zero(\$234\); default_zero(\$v1565\); default_zero(a); 
          default_zero(\$1228\); default_zero(\$861\); 
          default_zero(\$v3795\); default_zero(\$v3124\); 
          default_zero(\$v2549\); default_zero(\$v1982\); 
          default_zero(\$272\); default_zero(\$v2949\); 
          default_zero(\$v3388\); default_zero(\$v16_lock\); 
          default_zero(\$1195_i\); default_zero(\$739_lock\); 
          default_zero(\$v3272\); default_zero(\$v2286\); 
          default_zero(\$v4211\); default_zero(\$1417\); 
          default_zero(\$658\); default_zero(\$v2125\); 
          default_zero(\$v2302\); default_zero(\$436\); 
          default_zero(\$597_lock\); default_zero(\$689\); 
          default_zero(\$v1534\); default_zero(\$890\); 
          default_zero(\$874_lock\); default_zero(\$1562\); 
          default_zero(\$v1597\); default_zero(\$v3891\); 
          default_zero(\$452\); default_zero(\$444\); default_zero(\$v1815\); 
          default_zero(\$1220\); default_zero(\$1628\); 
          default_zero(\$571_lock\); default_zero(\$v3652\); 
          default_zero(\$705_lock\); default_zero(\$1178\); 
          default_zero(\$759\); default_zero(\$v2019\); default_zero(\$418\); 
          default_zero(\$v3113\); default_zero(\$653\); 
          default_zero(\$1084\); default_zero(\$v1702\); 
          default_zero(\$1390_lock\); default_zero(\$1119\); 
          default_zero(\$229\); default_zero(\$v2348\); 
          default_zero(\$1500\); default_zero(\$1080\); default_zero(\$500\); 
          default_zero(\$v3386\); default_zero(\$205\); 
          default_zero(\$1558\); default_zero(\$494\); 
          default_zero(\$v3141\); default_zero(\$1203_lock\); 
          default_zero(\$1529\); default_zero(\$v3370\); 
          default_zero(\$1618\); default_zero(\$v4079\); 
          default_zero(\$750\); default_zero(\$v30\); default_zero(\$v3705\); 
          default_zero(\$472\); default_zero(\$401_i\); 
          default_zero(\$v3120\); default_zero(\$v4206\); 
          default_zero(\$382\); default_zero(sp); default_zero(\$907\); 
          default_zero(\$1243\); default_zero(\$v2825\); 
          default_zero(\$981\); default_zero(\$v3234\); 
          default_zero(\$v2357\); default_zero(\$v2744\); 
          default_zero(\$v1473\); default_zero(\$v3495\); 
          default_zero(\$984_lock\); default_zero(\$v3431\); 
          default_zero(\$v3104\); default_zero(\$1354\); 
          default_zero(\$1287\); default_zero(\$v2226\); 
          default_zero(\$384\); default_zero(\$464_i\); 
          default_zero(\$1407\); default_zero(\$1468\); 
          default_zero(\$1339\); default_zero(\$1263_i\); 
          default_zero(\$1193\); default_zero(\$163\); default_zero(\$827\); 
          default_zero(\$v1983\); default_zero(\$v2865\); 
          default_zero(\$228\); default_zero(\$1174\); default_zero(\$482\); 
          default_zero(\$v2388\); default_zero(\$v3369\); 
          default_zero(\$v3433\); default_zero(\$v2599\); 
          default_zero(\$v3804\); default_zero(\$v1502\); 
          default_zero(\$1408\); default_zero(\$687_lock\); 
          default_zero(\$506_lock\); default_zero(\$1492_lock\); 
          default_zero(\$v1499\); default_zero(\$v3949\); 
          default_zero(\$v100\); default_zero(\$1255\); 
          default_zero(\$1180\); default_zero(\$1286\); 
          default_zero(\$947_lock\); default_zero(\$751\); 
          default_zero(\$v2829\); default_zero(\$364\); 
          default_zero(\$289_lock\); default_zero(\$v3310\); 
          default_zero(\$445\); default_zero(\$v3956\); default_zero(ib); 
          default_zero(\$v1756\); default_zero(\$v2354\); 
          default_zero(\$1357\); default_zero(\$486\); 
          default_zero(\$1074_x\); default_zero(\$v3745\); 
          default_zero(\$327\); default_zero(\$v1570\); 
          default_zero(\$1608\); default_zero(\$v1820\); 
          default_zero(\$v1624\); default_zero(\$1015\); 
          default_zero(\$1399\); default_zero(\$1138_lock\); 
          default_zero(\$1328_lock\); default_zero(\$v2179\); 
          default_zero(\$v1552\); default_zero(\$1031\); 
          default_zero(\$1010\); default_zero(\$v1956\); 
          default_zero(\$v3095\); default_zero(\$314\); 
          default_zero(\$v1484\); default_zero(\$795\); default_zero(\$544\); 
          default_zero(\$217\); default_zero(\$v2631\); 
          default_zero(\$1055\); default_zero(\$1248_lock\); 
          default_zero(\$v1529\); default_zero(\$v3669\); 
          default_zero(\$v32\); default_zero(\$178_lock\); 
          default_zero(\$v4084\); default_zero(\$705\); 
          default_zero(\$954_lock\); default_zero(\$v2996\); 
          default_zero(\$1462\); default_zero(\$v3437\); 
          default_zero(\$364_lock\); default_zero(\$850\); 
          default_zero(\$647\); default_zero(\$v36\); default_zero(\$v3597\); 
          default_zero(\$220_lock\); default_zero(\$81_i\); 
          default_zero(\$474\); default_zero(\$v3382\); 
          default_zero(\$v2198\); default_zero(\$617_lock\); 
          default_zero(\$982\); default_zero(\$v2749\); 
          default_zero(\$v3068\); default_zero(\$1348_lock\); 
          default_zero(\$1073\); default_zero(\$v3337\); 
          default_zero(\$v3798\); default_zero(\$v2330\); 
          default_zero(\$v3984\); default_zero(\$572\); default_zero(\$556\); 
          default_zero(\$v2262\); default_zero(\$1675_lock\); 
          default_zero(\$704\); default_zero(\$707_lock\); 
          default_zero(\$546\); default_zero(\$v2915\); 
          default_zero(\$1443\); default_zero(\$778\); default_zero(\$200\); 
          default_zero(\$1268_lock\); default_zero(\$164\); 
          default_zero(\$743_lock\); default_zero(\$69_x\); 
          default_zero(\$v2432\); default_zero(\$1448\); 
          default_zero(\$1168\); default_zero(\$v2618\); 
          default_zero(\$1069_lock\); default_zero(\$941\); 
          default_zero(\$255_lock\); default_zero(\$v3149\); 
          default_zero(\$1124_lock\); default_zero(\$177\); 
          default_zero(\$560\); default_zero(\$493\); default_zero(\$v2771\); 
          default_zero(\$732\); default_zero(\$618\); default_zero(\$1375\); 
          default_zero(\$254\); default_zero(\$v4029\); 
          default_zero(\$v1733\); default_zero(\$1022\); 
          default_zero(\$673_lock\); default_zero(\$v3638\); 
          default_zero(\$1125_result\); default_zero(\$1445\); 
          default_zero(\$566\); default_zero(\$v4034\); 
          default_zero(\$747_x\); default_zero(\$v2329\); 
          default_zero(\$435\); default_zero(\$v22\); default_zero(\$v2613\); 
          default_zero(\$1095\); default_zero(\$1262\); 
          default_zero(\$v2943\); default_zero(\$v3800\); 
          default_zero(\$591\); default_zero(\$v2408\); 
          default_zero(\$1557\); default_zero(\$598\); 
          default_zero(\$v2428\); default_zero(\$v3267\); 
          default_zero(\$v3822\); default_zero(\$v3461\); 
          default_zero(\$v1472\); default_zero(\$1267_lock\); 
          default_zero(\$1655\); default_zero(\$950_i\); 
          default_zero(\$v2419\); default_zero(\$v4193\); 
          default_zero(\$v4054\); default_zero(\$v1588\); 
          default_zero(\$1097\); default_zero(\$1482\); 
          default_zero(\$v3257\); default_zero(\$v3250\); 
          default_zero(\$1257\); default_zero(\$281\); 
          default_zero(\$1356_lock\); default_zero(\$1269\); 
          default_zero(\$v1618\); default_zero(\$v19_lock\); 
          default_zero(\$v3488\); default_zero(\$v3699\); 
          default_zero(\$v3831\); default_zero(\$856_x\); 
          default_zero(\$700\); default_zero(\$v2506\); 
          default_zero(\$1205\); default_zero(\$v2228\); 
          default_zero(\$v2600\); default_zero(\$968\); 
          default_zero(\$v2504\); default_zero(\$873_lock\); 
          default_zero(\$480\); default_zero(\$61_y\); 
          default_zero(\$v3965\); default_zero(\$v4125\); 
          default_zero(\$838_lock\); default_zero(\$v2418\); 
          default_zero(\$268\); default_zero(\$v3547\); 
          default_zero(\$352_lock\); default_zero(\$v3256\); 
          default_zero(\$607\); default_zero(\$v2036\); 
          default_zero(\$v3154\); default_zero(\$1045\); 
          default_zero(\$v2280\); default_zero(\$v2211\); 
          default_zero(\$v2204\); default_zero(\$v106\); 
          default_zero(\$v4116\); default_zero(\$v3897\); 
          default_zero(\$606\); default_zero(\$v3614\); 
          default_zero(\$1571_lock\); default_zero(\$326\); 
          default_zero(\$1395_lock\); default_zero(\$v3063\); 
          default_zero(\$668\); default_zero(\$476\); default_zero(\$v3884\); 
          default_zero(\$52_x\); default_zero(\$959_lock\); 
          default_zero(\$1530\); default_zero(\$56_y\); default_zero(\$419\); 
          default_zero(\$v1524\); default_zero(\$643\); default_zero(\$588\); 
          default_zero(\$v3392\); default_zero(\$v2042\); 
          default_zero(\$1237\); default_zero(\$v1606\); 
          default_zero(\$v1864\); default_zero(\$852_i\); 
          default_zero(\$v4146\); default_zero(\$v2096\); 
          default_zero(\$757\); default_zero(\$687\); default_zero(\$727\); 
          default_zero(\$329_lock\); default_zero(\$v2681\); 
          default_zero(\$1649\); default_zero(\$v3790\); 
          default_zero(\$59_tos\); default_zero(\$604_lock\); 
          default_zero(\$v93\); default_zero(\$v95\); default_zero(\$v1859\); 
          default_zero(\$571\); default_zero(\$437\); default_zero(\$349\); 
          default_zero(\$1281\); default_zero(\$714\); 
          default_zero(\$v3429\); default_zero(\$v38\); 
          default_zero(\$1569_lock\); default_zero(\$74_result_after_f\); 
          default_zero(\$868\); default_zero(\$810\); default_zero(\$v2676\); 
          default_zero(\$928\); default_zero(\$309_lock\); 
          default_zero(\$v3604\); default_zero(\$v2089\); 
          default_zero(\$v4121\); default_zero(\$301_lock\); 
          default_zero(\$v2248\); default_zero(\$v3091\); 
          default_zero(\$562_i\); default_zero(\$1601\); 
          default_zero(\$1497\); default_zero(\$v3126\); 
          default_zero(\$v2991\); default_zero(\$v1575\); 
          default_zero(\$1426\); default_zero(\$v3244\); 
          default_zero(\$1670\); default_zero(\$v3629\); 
          default_zero(\$206\); default_zero(\$970\); default_zero(\$v1684\); 
          default_zero(\$v3483\); default_zero(\$389\); 
          default_zero(\$v3809\); default_zero(\$1368\); 
          default_zero(\$584\); default_zero(\$710_i\); 
          default_zero(\$1551_lock\); default_zero(\$602\); 
          default_zero(\$v1854\); default_zero(\$960_x\); 
          default_zero(\$v4148\); default_zero(\$v3768\); 
          default_zero(\$1474\); default_zero(\$v4053\); 
          default_zero(\$v2480\); default_zero(\$519_lock\); 
          default_zero(\$1393\); default_zero(\$v4097\); 
          default_zero(\$v2483\); default_zero(\$v3827\); 
          default_zero(\$v3046\); default_zero(\$1138\); 
          default_zero(\$v37\); default_zero(tb); default_zero(\$1516_lock\); 
          default_zero(\$v2684\); default_zero(\$786\); 
          default_zero(\$v2143\); default_zero(\$1316_i\); 
          default_zero(\$690\); default_zero(\$1629\); 
          default_zero(\$1324_lock\); default_zero(\$1192\); 
          default_zero(\$1144_i\); default_zero(\$1441\); 
          default_zero(\$1234_lock\); default_zero(\$v4236\); 
          default_zero(\$v1799\); default_zero(\$v4111\); 
          default_zero(\$579_lock\); default_zero(\$372\); 
          default_zero(\$383\); default_zero(\$v3720\); 
          default_zero(\$v3153\); default_zero(\$v3741\); 
          default_zero(\$v2175\); default_zero(\$1207\); 
          default_zero(\$1300\); default_zero(\$832_lock\); 
          default_zero(\$v2636\); default_zero(\$v3196\); 
          default_zero(\$509\); default_zero(\$v2798\); 
          default_zero(\$641_lock\); default_zero(\$v3592\); 
          default_zero(\$v2013\); default_zero(\$1382_lock\); 
          default_zero(\$v1511\); default_zero(\$v3950\); 
          default_zero(\$1304\); default_zero(\$1499_x\); 
          default_zero(\$659_lock\); default_zero(\$v2426\); 
          default_zero(\$v3920\); default_zero(\$v2430\); 
          default_zero(\$1619\); default_zero(\$290\); default_zero(\$66_y\); 
          default_zero(\$v2356\); default_zero(\$1137\); 
          default_zero(\$v2796\); default_zero(\$v3109\); 
          default_zero(\$227\); default_zero(\$v1747\); 
          default_zero(\$v2971\); default_zero(\$543\); 
          default_zero(\$v4197\); default_zero(\$v2728\); 
          default_zero(\$786_lock\); default_zero(\$v3415\); 
          default_zero(\$84_x\); default_zero(\$965_x\); 
          default_zero(\$1442_x\); default_zero(\$1415_lock\); 
          default_zero(\$281_lock\); default_zero(\$v2523\); 
          default_zero(\$912\); default_zero(\$v2780\); 
          default_zero(\$v2366\); default_zero(\$558_lock\); 
          default_zero(\$399\); default_zero(\$v1798\); 
          default_zero(\$1644_x\); default_zero(\$v3238\); 
          default_zero(\$v2704\); default_zero(\$1097_lock\); 
          default_zero(\$1207_lock\); default_zero(\$1609\); 
          default_zero(\$505\); default_zero(\$v1731\); default_zero(\$162\); 
          default_zero(\$v2165\); default_zero(\$214_lock\); 
          default_zero(\$1383_x\); default_zero(\$1501\); 
          default_zero(\$301\); default_zero(\$434\); 
          default_zero(\$1179_lock\); default_zero(\$v1520\); 
          default_zero(\$706\); default_zero(\$397_lock\); 
          default_zero(\$1551\); default_zero(\$1363\); 
          default_zero(\$v2866\); default_zero(\$532\); 
          default_zero(\$v1802\); default_zero(\$1569\); 
          default_zero(\$603_lock\); default_zero(\$v3599\); 
          default_zero(\$v3064\); default_zero(\$1473\); 
          default_zero(\$v2627\); default_zero(\$1586\); 
          default_zero(\$396_lock\); default_zero(\$999\); 
          default_zero(\$v1619\); default_zero(\$v2107\); 
          default_zero(\$v42\); default_zero(\$1090_lock\); 
          default_zero(\$438_lock\); default_zero(\$1289_lock\); 
          default_zero(\$811\); default_zero(\$v3991\); 
          default_zero(\$1105\); default_zero(\$545\); 
          default_zero(\$488_x\); default_zero(\$v2370\); 
          default_zero(\$v31\); default_zero(\$v111\); default_zero(\$1229\); 
          default_zero(\$67_z\); default_zero(\$443\); default_zero(\$1248\); 
          default_zero(\$182\); default_zero(\$v74\); default_zero(\$v91\); 
          default_zero(\$v3405\); default_zero(\$1043\); 
          default_zero(\$v3867\); default_zero(\$1166\); 
          default_zero(\$766_lock\); default_zero(\$708\); 
          default_zero(\$v1488\); default_zero(\$v4170\); 
          default_zero(\$895\); default_zero(\$v1743\); 
          default_zero(\$1525\); default_zero(\$1616\); default_zero(\$794\); 
          default_zero(\$427_result_after_f\); default_zero(\$1662\); 
          default_zero(\$504\); default_zero(\$904\); default_zero(\$644\); 
          default_zero(\$v3223\); default_zero(\$920\); default_zero(\$201\); 
          default_zero(\$287\); default_zero(\$v2285\); 
          default_zero(\$1406\); default_zero(\$v4055\); 
          default_zero(\$258\); default_zero(\$876\); default_zero(\$918\); 
          default_zero(\$1213_i\); default_zero(\$433_lock\); 
          default_zero(\$v3130\); default_zero(\$1452\); 
          default_zero(\$308\); default_zero(\$v2298\); 
          default_zero(\$1206\); default_zero(\$1004_lock\); 
          default_zero(\$428_i\); default_zero(\$v20\); 
          default_zero(\$1069\); default_zero(\$1637\); 
          default_zero(\$1075_i\); default_zero(\$v1506\); 
          default_zero(\$v2043\); default_zero(\$976_lock\); 
          default_zero(\$v1889\); default_zero(\$1217_x\); 
          default_zero(\$727_lock\); default_zero(\$664_i\); 
          default_zero(\$v3451\); default_zero(\$v2569\); 
          default_zero(\$v1629\); default_zero(\$v3125\); 
          default_zero(\$1578\); default_zero(\$v2533\); 
          default_zero(\$v2403\); default_zero(\$v3836\); 
          default_zero(\$173\); default_zero(\$1638\); 
          default_zero(\$v1800\); default_zero(\$1596\); 
          default_zero(rdy1455); default_zero(\$1518_lock\); 
          default_zero(\$1516\); default_zero(\$v2735\); 
          default_zero(\$v2842\); default_zero(\$1194_result\); 
          default_zero(\$947\); default_zero(\$1447\); 
          default_zero(\$1022_lock\); default_zero(\$779\); 
          default_zero(\$616\); default_zero(\$v3551\); 
          default_zero(\$v3319\); default_zero(\$1435_lock\); 
          default_zero(\$v3354\); default_zero(\$v1793\); 
          default_zero(\$1315\); default_zero(\$v2427\); 
          default_zero(\$v3472\); default_zero(\$v3251\); 
          default_zero(\$1678\); default_zero(\$v3750\); 
          default_zero(\$181\); default_zero(\$1592\); 
          default_zero(\$372_lock\); default_zero(\$v1984\); 
          default_zero(\$225\); default_zero(\$v2170\); 
          default_zero(\$v1497\); default_zero(\$625_lock\); 
          default_zero(\$300\); default_zero(\$v1893\); 
          default_zero(\$640_lock\); default_zero(\$923\); 
          default_zero(\$v1865\); default_zero(result1454); 
          default_zero(\$460\); default_zero(\$691\); default_zero(\$1308\); 
          default_zero(\$792_lock\); default_zero(\$v1516\); 
          default_zero(\$1369\); default_zero(\$v2786\); 
          default_zero(\$256\); default_zero(\$1503\); 
          default_zero(\$v2266\); default_zero(\$v2431\); 
          default_zero(\$v28\); default_zero(\$719\); default_zero(\$v3364\); 
          default_zero(\$v3906\); default_zero(\$v3500\); 
          default_zero(\$733_lock\); default_zero(\$v1505\); 
          default_zero(\$v4184\); default_zero(\$v3754\); 
          default_zero(\$v1993\); default_zero(\$1676\); 
          default_zero(\$v1483\); default_zero(\$453\); 
          default_zero(\$v2787\); default_zero(\$1413_lock\); 
          default_zero(\$1555\); default_zero(\$645\); default_zero(\$1519\); 
          default_zero(\$v2018\); default_zero(\$424_lock\); 
          default_zero(\$385\); default_zero(\$199\); default_zero(\$v3774\); 
          default_zero(\$v1869\); default_zero(\$317_y\); 
          default_zero(\$1458\); default_zero(\$648\); 
          default_zero(\$v3730\); default_zero(\$1037\); 
          default_zero(\$660_lock\); default_zero(\$v4190\); 
          default_zero(\$v2792\); default_zero(\$738_lock\); 
          default_zero(\$1553\); default_zero(\$v3996\); 
          default_zero(\$v3059\); default_zero(\$586_x\); 
          default_zero(\$v2119\); default_zero(\$405\); 
          default_zero(\$1158\); default_zero(\$v3442\); 
          default_zero(\$1142_lock\); default_zero(\$v3992\); 
          default_zero(\$v2425\); default_zero(\$v2044\); 
          default_zero(\$991\); default_zero(\$v3907\); 
          default_zero(\$v2275\); default_zero(\$1056_lock\); 
          default_zero(\$v2034\); default_zero(\$620\); default_zero(\$824\); 
          default_zero(\$1473_lock\); default_zero(\$1340\); 
          default_zero(\$v3082\); default_zero(\$1005\); 
          default_zero(\$1584\); default_zero(\$1261\); 
          default_zero(\$v3317\); default_zero(\$v3943\); 
          default_zero(\$1333_i\); default_zero(\$v4011\); 
          default_zero(\$448\); default_zero(\$v3014\); 
          default_zero(\$v2116\); default_zero(\$1689\); 
          default_zero(\$319_i\); default_zero(\$v3799\); 
          default_zero(\$v3023\); default_zero(\$v2401\); 
          default_zero(\$764\); default_zero(\$v2611\); default_zero(\$587\); 
          default_zero(\$v1957\); default_zero(\$499\); 
          default_zero(\$135_i\); default_zero(\$v1841\); 
          default_zero(\$v1687\); default_zero(\$481\); 
          default_zero(\$v3137\); default_zero(\$v3490\); 
          default_zero(\$v2219\); default_zero(\$v1653\); 
          default_zero(\$v3383\); default_zero(\$985\); default_zero(\$172\); 
          default_zero(\$302\); default_zero(\$v1683\); 
          default_zero(\$v2560\); default_zero(\$v1688\); 
          default_zero(\$v2793\); default_zero(\$v3980\); 
          default_zero(\$1389_lock\); default_zero(\$936\); 
          default_zero(\$1096\); default_zero(\$1624\); 
          default_zero(\$1609_lock\); default_zero(\$255\); 
          default_zero(\$v3187\); default_zero(\$v1912\); 
          default_zero(\$1382\); default_zero(\$1056\); 
          default_zero(\$v2307\); default_zero(\$v3301\); 
          default_zero(\$1460_lock\); default_zero(\$v3974\); 
          default_zero(\$v120\); default_zero(\$v2852\); 
          default_zero(\$1187\); default_zero(\$v2662\); 
          default_zero(\$v2902\); default_zero(\$210_i\); 
          default_zero(\$933\); default_zero(\$1032\); 
          default_zero(\$1050_lock\); default_zero(\$526\); 
          default_zero(\$1400\); default_zero(\$693\); default_zero(\$1247\); 
          default_zero(\$1320_lock\); default_zero(\$1169\); 
          default_zero(\$v2492\); default_zero(\$1401\); 
          default_zero(\$v75\); default_zero(\$v3430\); 
          default_zero(\$1359_i\); default_zero(\$v2465\); 
          default_zero(\$v2045\); default_zero(\$v3854\); 
          default_zero(\$v3020\); default_zero(\$v3593\); 
          default_zero(\$659\); default_zero(\$35_a\); default_zero(\$1149\); 
          default_zero(\$323_lock\); default_zero(\$1117\); 
          default_zero(\$v3164\); default_zero(\$v2685\); 
          default_zero(\$1629_lock\); default_zero(\$1051\); 
          default_zero(\$v2802\); default_zero(\$462\); 
          default_zero(\$v3387\); default_zero(\$765_lock\); 
          default_zero(\$243_lock\); default_zero(\$v3492\); 
          default_zero(\$438\); default_zero(\$v4224\); 
          default_zero(\$v1811\); default_zero(\$v2410\); 
          default_zero(\$v4165\); default_zero(\$v1770\); 
          default_zero(\$758\); default_zero(\$v3961\); 
          default_zero(\$1148_x\); default_zero(\$v2663\); 
          default_zero(\$810_lock\); default_zero(\$v1852\); 
          default_zero(\$1598_x\); default_zero(\$v3990\); 
          default_zero(\$v2703\); default_zero(\$722\); 
          default_zero(\$v2929\); default_zero(\$v4122\); 
          default_zero(\$v3618\); default_zero(\$v2654\); 
          default_zero(\$840_y\); default_zero(\$v1678\); 
          default_zero(\$v4143\); default_zero(\$v1761\); 
          default_zero(\$v3159\); default_zero(\$v3291\); 
          default_zero(\$1517\); default_zero(\$v2537\); 
          default_zero(\$v3214\); default_zero(\$681\); default_zero(\$458\); 
          default_zero(\$1310\); default_zero(\$983\); 
          default_zero(\$v2659\); default_zero(\$1028\); 
          default_zero(\$681_lock\); default_zero(\$1428\); 
          default_zero(\$597\); default_zero(\$1165_lock\); 
          default_zero(\$1290\); default_zero(\$v3777\); 
          default_zero(\$v16\); default_zero(\$1664\); default_zero(\$423\); 
          default_zero(\$1249\); default_zero(\$1011_x\); 
          default_zero(\$v3543\); default_zero(\$v3776\); 
          default_zero(\$v2152\); default_zero(\$v3494\); 
          default_zero(\$v3087\); default_zero(\$324_lock\); 
          default_zero(\$v2856\); default_zero(\$v3619\); 
          default_zero(\$v2815\); default_zero(\$207_x\); 
          default_zero(\$v3169\); default_zero(\$1444\); 
          default_zero(\$v27_lock\); default_zero(\$1222\); 
          default_zero(\$v2234\); default_zero(\$1073_lock\); 
          default_zero(\$v2967\); default_zero(\$1337_x\); 
          default_zero(\$v1654\); default_zero(\$v4147\); 
          default_zero(\$v1548\); default_zero(\$v73\); 
          default_zero(\$996_lock\); default_zero(\$53_y\); 
          default_zero(\$1179\); default_zero(\$1033_i\); 
          default_zero(\$v2843\); default_zero(\$242\); 
          default_zero(\$v3666\); default_zero(\$1150\); 
          default_zero(\$v1707\); default_zero(\$v3465\); 
          default_zero(\$v3625\); default_zero(\$v3970\); 
          default_zero(\$v2622\); default_zero(\$1143_x\); 
          default_zero(\$v1677\); default_zero(\$1256_lock\); 
          default_zero(\$v3410\); default_zero(\$32_a\); 
          default_zero(\$v2130\); default_zero(\$v2601\); 
          default_zero(\$728\); default_zero(\$796\); default_zero(\$336\); 
          default_zero(\$282\); default_zero(\$v3365\); 
          default_zero(\$v1711\); default_zero(\$v2978\); 
          default_zero(\$191\); default_zero(\$1301\); default_zero(\$269\); 
          default_zero(\$851_x\); default_zero(\$1459\); 
          default_zero(\$390_lock\); default_zero(\$v3634\); 
          default_zero(\$v2727\); default_zero(\$1013\); 
          default_zero(\$875_lock\); default_zero(\$1647\); 
          default_zero(\$520\); default_zero(\$460_lock\); 
          default_zero(\$373\); default_zero(\$557_lock\); 
          default_zero(\$1510\); default_zero(\$208_y\); 
          default_zero(\$v3191\); default_zero(\$171\); 
          default_zero(\$1414_lock\); default_zero(\$v4089\); 
          default_zero(\$803\); default_zero(\$522\); 
          default_zero(\$1042_lock\); default_zero(\$1349\); 
          default_zero(\$v3501\); default_zero(\$v3000\); 
          default_zero(\$487_lock\); default_zero(\$55_x\); 
          default_zero(\$v1732\); default_zero(\$350\); 
          default_zero(\$v1860\); default_zero(\$v3841\); 
          default_zero(\$v1914\); default_zero(\$1568\); 
          default_zero(\$1453_lock\); default_zero(\$966\); 
          default_zero(\$v2740\); default_zero(\$v2002\); 
          default_zero(\$903\); default_zero(\$1096_lock\); 
          default_zero(\$v4202\); default_zero(\$v4123\); 
          default_zero(\$398_lock\); default_zero(\$995\); 
          default_zero(\$1436\); default_zero(\$v3283\); 
          default_zero(\$v3218\); default_zero(\$377\); 
          default_zero(\$v4166\); default_zero(\$1029\); 
          default_zero(\$v1471\); default_zero(\$1338\); 
          default_zero(\$264\); default_zero(\$v3546\); default_zero(\$748\); 
          default_zero(\$v2451\); default_zero(\$631_lock\); 
          default_zero(\$v2950\); default_zero(\$v3511\); 
          default_zero(\$418_lock\); default_zero(\$720\); 
          default_zero(\$1309_lock\); default_zero(\$673\); 
          default_zero(\$v1573\); default_zero(\$v2098\); 
          default_zero(\$1199_lock\); default_zero(\$652\); 
          default_zero(\$1170_i\); default_zero(\$v1988\); 
          default_zero(\$v2579\); default_zero(\$v3670\); 
          default_zero(\$1165\); default_zero(pos); default_zero(\$v3565\); 
          default_zero(\$v2053\); default_zero(\$367\); 
          default_zero(\$1549_lock\); default_zero(\$1354_lock\); 
          default_zero(\$v2729\); default_zero(\$v35\); 
          default_zero(\$1563_lock\); default_zero(\$1414\); 
          default_zero(\$1081\); default_zero(\$304\); 
          default_zero(\$v3524\); default_zero(\$1091\); 
          default_zero(\$1675\); default_zero(\$961_i\); 
          default_zero(\$73_result\); default_zero(\$1212_x\); 
          default_zero(\$v2589\); default_zero(\$1498_lock\); 
          default_zero(\$v3642\); default_zero(\$514\); 
          default_zero(\$v1467\); default_zero(\$527\); default_zero(\$672\); 
          default_zero(\$v2635\); default_zero(\$v1616\); 
          default_zero(\$v2870\); default_zero(\$1454\); 
          default_zero(\$v3661\); default_zero(\$v4030\); 
          default_zero(\$v1706\); default_zero(\$v3544\); 
          default_zero(\$798\); default_zero(\$v3902\); 
          default_zero(\$1689_lock\); default_zero(\$v2417\); 
          default_zero(\$686\); default_zero(\$608_i\); default_zero(\$676\); 
          default_zero(\$1650\); default_zero(\$v1997\); 
          default_zero(\$1550_lock\); default_zero(\$579\); 
          default_zero(\$v3227\); default_zero(\$v3896\); 
          default_zero(\$585_lock\); default_zero(\$906\); 
          default_zero(\$1050\); default_zero(\$653_lock\); 
          default_zero(\$65_x\); default_zero(\$1269_lock\); 
          default_zero(\$624\); default_zero(\$v3951\); 
          default_zero(\$v3381\); default_zero(\$1688\); 
          default_zero(\$v2120\); default_zero(\$1418_i\); 
          default_zero(\$275\); default_zero(\$v2897\); 
          default_zero(\$328_lock\); default_zero(\$161_x\); 
          default_zero(\$v2017\); default_zero(\$719_lock\); 
          default_zero(\$v1875\); default_zero(\$v3178\); 
          default_zero(\$76_result\); default_zero(\$674\); 
          default_zero(\$v3352\); default_zero(\$v3916\); 
          default_zero(\$896\); default_zero(\$1003\); default_zero(\$781\); 
          default_zero(\$219_lock\); default_zero(\$1142\); 
          default_zero(\$v3376\); default_zero(\$1061_lock\); 
          default_zero(\$1275\); default_zero(\$v3205\); 
          default_zero(\$v1939\); default_zero(\$355_i\); 
          default_zero(\$1272\); default_zero(\$1065_lock\); 
          default_zero(\$v2261\); default_zero(\$v2334\); 
          default_zero(\$1460\); default_zero(\$v2218\); 
          default_zero(\$v2066\); default_zero(ta); 
          default_zero(\$437_lock\); default_zero(\$574\); 
          default_zero(\$400\); default_zero(\$v2781\); 
          default_zero(\$1238\); default_zero(\$1517_lock\); 
          default_zero(\$v3736\); default_zero(\$241_lock\); 
          default_zero(\$v40\); default_zero(\$v2505\); 
          default_zero(\$v1784\); default_zero(\$v3424\); 
          default_zero(\$1570\); default_zero(\$v1633\); 
          default_zero(\$v3715\); default_zero(\$v3021\); 
          default_zero(\$v1525\); default_zero(\$542\); default_zero(\$777\); 
          default_zero(\$v2139\); default_zero(\$v2791\); 
          default_zero(\$v3773\); default_zero(\$v17\); 
          default_zero(\$1042\); default_zero(\$1066\); 
          default_zero(\$v3721\); default_zero(\$787\); 
          default_zero(\$v1489\); default_zero(\$1367\); 
          default_zero(\$v2820\); default_zero(\$v2769\); 
          default_zero(\$v1620\); default_zero(\$592\); 
          default_zero(\$v1961\); default_zero(\$v3587\); 
          default_zero(\$v3613\); default_zero(\$823\); default_zero(\$310\); 
          default_zero(\$v3520\); default_zero(\$642_x\); 
          default_zero(\$v2775\); default_zero(\$1407_lock\); 
          default_zero(\$1204\); default_zero(\$785\); default_zero(\$1683\); 
          default_zero(\$631\); default_zero(\$180_lock\); 
          default_zero(\$v2271\); default_zero(\$v1806\); 
          default_zero(\$v3842\); default_zero(\$1487_lock\); 
          default_zero(\$v2487\); default_zero(\$533\); 
          default_zero(\$v2909\); default_zero(\$v1659\); default_zero(pc); 
          default_zero(\$1239_i\); default_zero(\$765\); 
          default_zero(\$1645\); default_zero(\$v2035\); 
          default_zero(\$1017\); default_zero(\$1502\); 
          default_zero(\$v1655\); default_zero(\$1554\); 
          default_zero(\$236\); default_zero(\$1663_lock\); 
          default_zero(\$604\); default_zero(result); default_zero(\$v1734\); 
          default_zero(\$v3843\); default_zero(\$1453\); 
          default_zero(\$934\); default_zero(\$1099\); default_zero(\$1358\); 
          default_zero(\$v1943\); default_zero(\$328\); 
          default_zero(\$1597\); default_zero(\$1110_lock\); 
          default_zero(\$1085\); default_zero(\$603\); 
          default_zero(\$v2385\); default_zero(\$v2134\); 
          default_zero(\$v2550\); default_zero(\$v3538\); 
          default_zero(\$v3036\); default_zero(\$550\); 
          default_zero(\$v2583\); default_zero(\$v3240\); 
          default_zero(\$335\); default_zero(\$v104\); 
          default_zero(\$1530_lock\); default_zero(\$v3667\); 
          default_zero(\$v4107\); default_zero(\$1603\); 
          default_zero(\$v3874\); default_zero(\$v3296\); 
          default_zero(\$1381\); default_zero(\$699_lock\); 
          default_zero(\$v1880\); default_zero(\$273\); 
          default_zero(\$v67_lock\); default_zero(\$447\); 
          default_zero(\$v2343\); default_zero(\$v2200\); 
          default_zero(\$949_y\); default_zero(\$v2390\); 
          default_zero(\$1521_i\); default_zero(\$1591_lock\); 
          default_zero(\$v2496\); default_zero(\$413\); 
          default_zero(\$1221\); default_zero(\$v3005\); 
          default_zero(\$1030_lock\); default_zero(\$v3255\); 
          default_zero(\$527_lock\); default_zero(\$1661\); 
          default_zero(\$v3598\); default_zero(\$v2995\); 
          default_zero(\$v2413\); default_zero(\$551\); 
          default_zero(\$v4098\); default_zero(\$v1981\); 
          default_zero(\$1012\); default_zero(\$v2288\); 
          default_zero(\$559_lock\); default_zero(\$v2289\); 
          default_zero(\$v1561\); default_zero(\$v2361\); 
          default_zero(\$v4025\); default_zero(\$v2722\); 
          default_zero(\$v2411\); default_zero(\$v3781\); 
          default_zero(\$490\); default_zero(\$561\); default_zero(\$v4048\); 
          default_zero(\$1187_lock\); default_zero(\$1661_lock\); 
          default_zero(\$743\); default_zero(\$v2884\); default_zero(\$380\); 
          default_zero(\$858\); default_zero(\$v1671\); default_zero(\$749\); 
          default_zero(\$v3278\); default_zero(\$v1689\); 
          default_zero(\$v76_lock\); default_zero(\$v2111\); 
          default_zero(\$v1498\); default_zero(\$v2391\); 
          default_zero(\$v2084\); default_zero(\$v3482\); 
          default_zero(\$v2959\); default_zero(\$1495\); 
          default_zero(\$v1788\); default_zero(\$v1861\); 
          default_zero(\$1531\); default_zero(\$v73_lock\); 
          default_zero(\$955_lock\); default_zero(\$824_lock\); 
          default_zero(\$1235\); default_zero(\$v2811\); 
          default_zero(\$v2409\); default_zero(\$v45_lock\); 
          default_zero(\$v3041\); default_zero(\$1642\); 
          default_zero(\$913_lock\); default_zero(\$768\); 
          default_zero(\$v39\); default_zero(\$v3496\); 
          default_zero(\$v2893\); default_zero(\$v3045\); 
          default_zero(\$1377\); default_zero(\$v2690\); 
          default_zero(\$315\); default_zero(\$1113\); 
          default_zero(\$793_x\); default_zero(\$v2287\); 
          default_zero(\$v3077\); default_zero(\$1079_x\); 
          default_zero(\$1511\); default_zero(\$1082\); 
          default_zero(\$v2244\); default_zero(\$1544_lock\); 
          default_zero(\$1602\); default_zero(\$v3323\); 
          default_zero(\$663\); default_zero(\$v3377\); default_zero(\$353\); 
          default_zero(\$v3692\); default_zero(\$1488_i\); 
          default_zero(\$378\); default_zero(\$v2429\); default_zero(\$959\); 
          default_zero(\$v4189\); default_zero(\$1464_i\); 
          default_zero(\$1537\); default_zero(\$71_result_after_f\); 
          default_zero(\$v4102\); default_zero(\$v3142\); 
          default_zero(\$882\); default_zero(\$v2048\); default_zero(\$325\); 
          default_zero(\$v2148\); default_zero(\$v2212\); 
          default_zero(\$558\); default_zero(\$v1752\); 
          default_zero(\$769_i\); default_zero(\$v3305\); 
          default_zero(\$v96\); default_zero(\$v1549\); 
          default_zero(\$442_x\); default_zero(\$v2041\); 
          default_zero(\$v2239\); default_zero(\$v114\); 
          default_zero(\$v3506\); default_zero(\$v1952\); 
          default_zero(\$v4179\); default_zero(\$343\); 
          default_zero(\$1397\); default_zero(\$v2402\); 
          default_zero(\$1582\); default_zero(\$v2166\); 
          default_zero(\$v1584\); default_zero(\$1110\); 
          default_zero(\$1539\); default_zero(\$1476\); 
          default_zero(\$v2911\); default_zero(\$1660\); 
          default_zero(\$v89\); default_zero(\$1648\); 
          default_zero(\$v2555\); default_zero(\$172_lock\); 
          default_zero(\$1563\); default_zero(\$v3576\); 
          default_zero(\$1314\); default_zero(\$1656\); 
          default_zero(\$v1593\); default_zero(\$v3032\); 
          default_zero(\$v3580\); default_zero(\$v2242\); 
          default_zero(\$287_lock\); default_zero(\$v4000\); 
          default_zero(\$975\); default_zero(\$1282\); 
          default_zero(\$v2528\); default_zero(\$v78_lock\); 
          default_zero(\$1009\); default_zero(\$v2982\); 
          default_zero(\$v2023\); default_zero(\$379_x\); 
          default_zero(\$v4057\); default_zero(\$v2816\); 
          default_zero(\$226\); default_zero(\$187\); default_zero(\$v2939\); 
          default_zero(\$v1507\); default_zero(\$1332_x\); 
          default_zero(\$1211_lock\); default_zero(\$v2195\); 
          default_zero(\$v3136\); default_zero(\$v3533\); 
          default_zero(\$v2960\); default_zero(\$v3515\); 
          default_zero(\$838\); default_zero(\$682\); default_zero(\$541\); 
          default_zero(\$v2163\); default_zero(\$v2094\); 
          default_zero(\$v1866\); default_zero(\$1446\); 
          default_zero(\$v3716\); default_zero(\$351\); default_zero(\$245\); 
          default_zero(\$200_lock\); default_zero(\$v4129\); 
          default_zero(\$v2840\); default_zero(\$v2102\); 
          default_zero(\$v2257\); default_zero(\$1498\); 
          default_zero(\$v3588\); default_zero(\$1493_lock\); 
          default_zero(\$v3358\); default_zero(\$v2395\); 
          default_zero(\$241\); default_zero(\$v3088\); 
          default_zero(\$v4016\); default_zero(\$1614\); 
          default_zero(\$1481_lock\); default_zero(\$390\); 
          default_zero(\$82_i\); default_zero(\$932\); 
          default_zero(\$v4021\); default_zero(\$1682\); 
          default_zero(\$1427\); default_zero(ia); default_zero(\$424\); 
          default_zero(\$694\); default_zero(\$914\); default_zero(\$v2551\); 
          default_zero(\$886\); default_zero(\$v1920\); 
          default_zero(\$v4192\); default_zero(\$v2606\); 
          default_zero(\$1233\); default_zero(\$v3924\); 
          default_zero(\$1505\); default_zero(\$v2661\); 
          default_zero(\$v2708\); default_zero(\$192\); 
          default_zero(\$1376\); default_zero(\$1126_i\); 
          default_zero(\$v1720\); default_zero(\$179\); 
          default_zero(\$209_result_after_f\); default_zero(\$v3201\); 
          default_zero(\$v2311\); default_zero(\$v2046\); 
          default_zero(\$1193_lock\); default_zero(\$758_lock\); 
          default_zero(\$873\); default_zero(\$v1642\); 
          default_zero(\$v2645\); default_zero(\$v2924\); 
          default_zero(\$v2807\); default_zero(\$v2797\); 
          default_zero(\$v23\); default_zero(\$982_lock\); 
          default_zero(\$718\); default_zero(stbl); default_zero(\$1152\); 
          default_zero(\$551_lock\); default_zero(\$557\); 
          default_zero(\$902_x\); default_zero(\$v2987\); 
          default_zero(\$v2847\); default_zero(\$v4010\); 
          default_zero(\$976\); default_zero(\$v2510\); 
          default_zero(\$v2841\); default_zero(\$235_lock\); 
          default_zero(\$1288_lock\); default_zero(\$1273\); 
          default_zero(\$654\); default_zero(\$v3556\); default_zero(\$905\); 
          default_zero(\$276\); default_zero(\$v3009\); default_zero(\$381\); 
          default_zero(\$v2051\); default_zero(\$920_lock\); 
          default_zero(\$986\); default_zero(\$v2162\); 
          default_zero(\$1023\); default_zero(\$1441_lock\); 
          default_zero(\$v45\); default_zero(\$v4161\); 
          default_zero(\$473_lock\); default_zero(\$v4078\); 
          default_zero(\$v2216\); default_zero(\$v2316\); 
          default_zero(\$v31_lock\); default_zero(\$942\); 
          default_zero(\$506\); default_zero(\$941_lock\); 
          default_zero(\$933_lock\); default_zero(\$908\); 
          default_zero(\$1662_lock\); default_zero(\$v3481\); 
          default_zero(\$1057_i\); default_zero(\$v3493\); 
          default_zero(\$1533\); default_zero(\$924_i\); 
          default_zero(\$v2447\); default_zero(\$167\); 
          default_zero(\$v2763\); default_zero(\$v44\); 
          default_zero(\$v2424\); default_zero(\$646\); default_zero(\$867\); 
          default_zero(\$1597_lock\); default_zero(\$1049\); 
          default_zero(\$v1579\); default_zero(\$137_i\); 
          default_zero(\$1256\); default_zero(\$v2861\); 
          default_zero(\$v1638\); default_zero(\$1228_lock\); 
          default_zero(\$271\); default_zero(\$v2548\); default_zero(\$v33\); 
          default_zero(\$v108\); default_zero(\$v4043\); 
          default_zero(\$v2973\); default_zero(\$1637_lock\); 
          default_zero(\$459_lock\); default_zero(\$1416\); 
          default_zero(\$v4240\); default_zero(\$940\); default_zero(\$v21\); 
          default_zero(\$v3027\); default_zero(\$v3890\); 
          default_zero(\$946\); default_zero(\$580\); default_zero(\$v3844\); 
          default_zero(\$v3100\); default_zero(\$v2375\); 
          default_zero(\$1276\); default_zero(\$v3209\); 
          default_zero(\$v3318\); default_zero(\$v1862\); 
          default_zero(\$v3732\); default_zero(\$v4134\); 
          default_zero(\$195\); default_zero(\$v1929\); 
          default_zero(\$1368_lock\); default_zero(\$866\); 
          default_zero(\$v1693\); default_zero(\$v3315\); 
          default_zero(\$1570_lock\); default_zero(\$578\); 
          default_zero(\$263\); default_zero(\$v2197\); 
          default_zero(\$v4075\); default_zero(\$v3160\); 
          default_zero(\$v2220\); default_zero(\$v2188\); 
          default_zero(\$1301_lock\); default_zero(\$1089\); 
          default_zero(\$971\); default_zero(\$1090\); 
          default_zero(\$v2238\); default_zero(\$v3239\); 
          default_zero(\$1348\); default_zero(\$v28_lock\); 
          default_zero(\$1599\); default_zero(\$v25\); default_zero(\$83_x\); 
          default_zero(\$1029_lock\); default_zero(\$333_x\); 
          default_zero(\$165\); default_zero(\$585\); default_zero(\$977\); 
          default_zero(\$492\); default_zero(\$v2199\); default_zero(\$612\); 
          default_zero(\$1655_lock\); default_zero(\$v3749\); 
          default_zero(\$230\); default_zero(\$841_i\); default_zero(\$468\); 
          default_zero(\$v79\); default_zero(\$v2164\); default_zero(\$463\); 
          default_zero(\$432_lock\); default_zero(\$1083\); 
          default_zero(\$v3273\); default_zero(\$850_lock\); 
          default_zero(\$1211\); default_zero(\$26_a\); 
          default_zero(\$1188\); default_zero(\$874\); default_zero(\$371\); 
          default_zero(\$v3262\); default_zero(\$996\); default_zero(\$832\); 
          default_zero(\$1186\); default_zero(\$v2933\); 
          default_zero(\$v4066\); default_zero(\$v3177\); 
          default_zero(\$280\); default_zero(\$812_lock\); 
          default_zero(\$v3050\); default_zero(\$v26\); 
          default_zero(\$v3813\); default_zero(\$318_result_after_f\); 
          default_zero(\$v1884\); default_zero(\$1041\); 
          default_zero(\$v3471\); default_zero(\$552\); default_zero(\$338\); 
          default_zero(\$1486\); default_zero(\$596\); 
          default_zero(\$v1980\); default_zero(\$605_lock\); 
          default_zero(\$v2047\); default_zero(\$v3477\); 
          default_zero(\$v2564\); default_zero(\$v3202\); 
          default_zero(\$v3786\); default_zero(\$1398\); 
          default_zero(\$639_lock\); default_zero(\$1014\); 
          default_zero(\$v1837\); default_zero(\$v3491\); 
          default_zero(\$1251\); default_zero(\$1182\); 
          default_zero(\$540_x\); default_zero(\$417\); 
          default_zero(\$v2217\); default_zero(\$1610\); 
          default_zero(\$v1779\); default_zero(\$v3679\); 
          default_zero(\$1234\); default_zero(\$1643\); 
          default_zero(\$1223\); default_zero(\$1227\); default_zero(\$v19\); 
          default_zero(\$v2412\); default_zero(\$1497_lock\); 
          default_zero(\$v1500\); default_zero(\$291\); 
          default_zero(\$v3575\); default_zero(\$837\); default_zero(\$831\); 
          default_zero(\$1292_i\); default_zero(\$v2121\); 
          default_zero(\$1646\); default_zero(\$1167_lock\); 
          default_zero(\$491\); default_zero(\$1459_lock\); 
          default_zero(\$1545_i\); default_zero(\$1291\); 
          default_zero(\$1151\); default_zero(\$206_lock\); 
          default_zero(\$v3090\); default_zero(\$833\); default_zero(\$967\); 
          default_zero(\$274\); default_zero(\$v2875\); 
          default_zero(\$1665\); default_zero(\$799\); 
          default_zero(\$633_y\); default_zero(\$v1682\); 
          default_zero(\$1100\); default_zero(\$498\); 
          default_zero(\$v2355\); default_zero(\$v1550\); 
          default_zero(\$1590\); default_zero(\$1028_lock\); 
          default_zero(\$922\); default_zero(\$v3925\); 
          default_zero(\$v2469\); default_zero(\$948_x\); 
          default_zero(\$v22_lock\); default_zero(\$v3489\); 
          default_zero(\$v3148\); default_zero(\$v27\); default_zero(\$894\); 
          default_zero(\$862\); default_zero(\$987_i\); 
          default_zero(\$v1755\); default_zero(\$1440\); 
          default_zero(\$v3569\); default_zero(\$391\); 
          default_zero(\$1591\); default_zero(\$v2006\); 
          default_zero(\$1068\); default_zero(\$1154\); 
          default_zero(\$316_x\); default_zero(\$v3703\); 
          default_zero(\$v2456\); default_zero(\$1643_lock\); 
          default_zero(\$v2442\); default_zero(\$v2029\); 
          default_zero(\$v3269\); default_zero(\$877\); 
          default_zero(\$v2433\); default_zero(\$v3624\); 
          default_zero(\$v2436\); default_zero(\$845_lock\); 
          default_zero(\$v2481\); default_zero(\$1016\); 
          default_zero(\$1219\); default_zero(\$v2237\); 
          default_zero(\$v55_lock\); default_zero(\$v3863\); 
          default_zero(\$v2353\); default_zero(\$1343\); 
          default_zero(\$v3348\); default_zero(\$1159\); 
          default_zero(\$698\); default_zero(\$v1490\); 
          default_zero(\$v3022\); default_zero(\$662\); 
          default_zero(\$1434\); default_zero(\$v3446\); 
          default_zero(\$v3455\); default_zero(\$v2612\); 
          default_zero(\$634_result\); default_zero(\$v4232\); 
          default_zero(\$v3529\); default_zero(\$410_lock\); 
          default_zero(\$397\); default_zero(b); default_zero(\$v2030\); 
          default_zero(\$v2387\); default_zero(\$v1847\); 
          default_zero(\$528\); default_zero(\$1101_i\); 
          default_zero(\$v2713\); default_zero(\$v3688\); 
          default_zero(\$v3643\); default_zero(\$1392\); 
          default_zero(\$v2883\); default_zero(\$224_x\); 
          default_zero(\$v4215\); default_zero(\$900\); default_zero(\$692\); 
          default_zero(\$v2640\); default_zero(\$1164\); 
          default_zero(\$v1848\); default_zero(\$1583\); 
          default_zero(\$1461_lock\); default_zero(\$v2547\); 
          default_zero(\$250\); default_zero(\$263_lock\); 
          default_zero(\$v3401\); default_zero(\$288_lock\); 
          default_zero(\$1376_lock\); default_zero(\$1136\); 
          default_zero(\$688_x\); default_zero(\$v3763\); 
          default_zero(\$1504\); default_zero(\$v3158\); 
          default_zero(\$246_i\); default_zero(\$454\); default_zero(\$216\); 
          default_zero(\$632_x\); default_zero(\$v117\); 
          default_zero(\$v1670\); default_zero(\$v3182\); 
          default_zero(\$v2519\); default_zero(\$1674\); 
          default_zero(\$1004\); default_zero(\$288\); 
          default_zero(\$v3709\); default_zero(\$v3341\); 
          default_zero(\$857\); default_zero(\$v3656\); 
          default_zero(\$v2972\); default_zero(\$v2138\); 
          default_zero(\$v2779\); default_zero(\$29_a\); 
          default_zero(\$v1824\); default_zero(\$v3328\); 
          default_zero(\$733\); default_zero(\$v3044\); 
          default_zero(\$1109\); default_zero(\$v3683\); 
          default_zero(\$v60_lock\); default_zero(\$v2437\); 
          default_zero(\$v1774\); default_zero(\$v78\); 
          default_zero(\$1355_lock\); default_zero(\$518\); 
          default_zero(\$339\); default_zero(\$1123\); 
          default_zero(\$v1666\); default_zero(\$v3948\); 
          default_zero(\$334\); default_zero(\$1515\); 
          default_zero(\$v1902\); default_zero(\$1402\); 
          default_zero(\$997\); default_zero(\$1574_i\); 
          default_zero(\$v3274\); default_zero(\$v1966\); 
          default_zero(\$v3775\); default_zero(\$v3316\); 
          default_zero(\$v4002\); default_zero(\$872\); 
          default_zero(\$1572\); default_zero(\$630\); 
          default_zero(\$v2057\); default_zero(\$1430\); 
          default_zero(\$797\); default_zero(\$1472\); 
          default_zero(\$v2955\); default_zero(\$1556\); 
          default_zero(\$1271\); default_zero(\$v1853\); 
          default_zero(\$v4124\); default_zero(\$1341\); 
          default_zero(\$v2907\); default_zero(\$v2479\); 
          default_zero(\$v2062\); default_zero(\$v1898\); 
          default_zero(\$425_x\); default_zero(\$v2695\); 
          default_zero(\$1270_x\); default_zero(\$v1538\); 
          default_zero(\$337\); default_zero(\$v1680\); 
          default_zero(\$v2864\); default_zero(\$811_lock\); 
          default_zero(\$v2253\); default_zero(\$v3406\); 
          default_zero(\$v3419\); default_zero(\$590\); 
          default_zero(\$315_lock\); default_zero(\$v3647\); 
          default_zero(\$v3608\); default_zero(\$v2233\); 
          default_zero(\$v3586\); default_zero(\$969\); default_zero(\$519\); 
          default_zero(\$v2590\); default_zero(\$v3911\); 
          default_zero(\$v94\); default_zero(\$v2243\); 
          default_zero(\$v1738\); default_zero(\$487\); 
          default_zero(\$v2196\); default_zero(\$269_lock\); 
          default_zero(\$v2293\); default_zero(\$v2839\); 
          default_zero(\$753\); default_zero(\$235\); default_zero(\$v3938\); 
          default_zero(\$v3704\); default_zero(\$v1730\); 
          default_zero(\$v2753\); default_zero(\$v3204\); 
          default_zero(\$1481\); default_zero(\$378_lock\); 
          default_zero(\$363\); default_zero(\$v3759\); 
          default_zero(\$901_lock\); default_zero(\$v1913\); 
          default_zero(\$v3497\); default_zero(\$v2616\); 
          default_zero(\$v1801\); default_zero(\$v41\); 
          default_zero(\$v2386\); default_zero(\$v3845\); 
          default_zero(\$v3818\); default_zero(\$v4001\); 
          default_zero(\$1287_lock\); default_zero(\$309\); 
          default_zero(\$461_lock\); default_zero(\$v2672\); 
          default_zero(\$v2438\); default_zero(\$1654\); 
          default_zero(\$767\); default_zero(\$v3668\); 
          default_zero(\$895_lock\); default_zero(\$296\); 
          default_zero(\$v3623\); default_zero(\$v2321\); 
          default_zero(\$773\); default_zero(\$218\); default_zero(\$791\); 
          default_zero(\$726\); default_zero(\$v3895\); 
          default_zero(\$v2888\); default_zero(\$v2951\); 
          default_zero(\$351_lock\); default_zero(\$v1460\); 
          default_zero(\$365\); default_zero(\$v3731\); 
          default_zero(\$v1679\); default_zero(\$1309\); 
          default_zero(\$344_lock\); default_zero(\$v3858\); 
          default_zero(\$1394_lock\); default_zero(\$v1501\); 
          default_zero(\$v80\); default_zero(\$v3268\); 
          default_zero(\$v3560\); default_zero(\$v1948\); 
          default_zero(\$1134_lock\); default_zero(\$v1496\); 
          default_zero(\$244\); default_zero(\$1422\); 
          default_zero(\$507_lock\); default_zero(\$v1870\); 
          default_zero(\$1630\); default_zero(\$706_lock\); 
          default_zero(\$v4157\); default_zero(\$270_x\); 
          default_zero(\$1021\); default_zero(\$v3089\); 
          default_zero(\$878_i\); default_zero(\$1098_lock\); 
          default_zero(\$v43_lock\); default_zero(\$v2770\); 
          default_zero(\$815_i\); default_zero(\$v3371\); 
          default_zero(\$v2184\); default_zero(\$1615_lock\); 
          default_zero(\$1342\); default_zero(\$1552_x\); 
          default_zero(\$v2407\); default_zero(\$v3073\); 
          default_zero(\$v1831\); default_zero(\$1604\); 
          default_zero(\$1636\); default_zero(\$v3905\); 
          default_zero(\$919_lock\); default_zero(\$v3929\); 
          default_zero(\$v2460\); default_zero(\$v2595\); 
          default_zero(\$v3203\); default_zero(\$813\); 
          default_zero(\$v2221\); default_zero(\$v3620\); 
          default_zero(\$921_lock\); default_zero(\$1600\); 
          default_zero(\$v1495\); default_zero(\$v2070\); 
          default_zero(\$v2717\); default_zero(\$262\); 
          default_zero(\$v2976\); default_zero(\$510_i\); 
          default_zero(\$v4061\); default_zero(\$v2667\); 
          default_zero(\$58_result\); default_zero(\$v2236\); 
          default_zero(\$v2455\); default_zero(\$1111\); 
          default_zero(\$v3952\); default_zero(\$1118_lock\); 
          default_zero(\$1583_lock\); default_zero(\$426_y\); 
          default_zero(\$v1907\); default_zero(\$1683_lock\); 
          default_zero(\$220\); default_zero(\$481_lock\); 
          default_zero(\$v2966\); default_zero(\$459\); 
          default_zero(\$v2759\); default_zero(\$660\); 
          default_zero(\$1617_lock\); default_zero(\$v2071\); 
          default_zero(\$v4039\); default_zero(\$v1937\); 
          default_zero(\$1435\); default_zero(\$395\); 
          default_zero(\$v2194\); default_zero(\$v1775\); 
          default_zero(\$901\); default_zero(\$v2591\); 
          default_zero(\$983_lock\); default_zero(\$v3879\); 
          default_zero(\$v1766\); default_zero(\$166\); default_zero(\$792\); 
          default_zero(\$396\); default_zero(\$v4093\); 
          default_zero(\$1274\); default_zero(\$v1477\); 
          default_zero(\$v4191\); default_zero(\$v1649\); 
          default_zero(\$v2389\); default_zero(\$v1665\); 
          default_zero(\$v1888\); default_zero(\$1510_lock\); 
          default_zero(\$v24\); default_zero(\$v3880\); 
          default_zero(\$1385_i\); default_zero(\$v1970\); 
          default_zero(\$v4070\); default_zero(\$1118\); 
          default_zero(\$v3155\); default_zero(\$v2977\); 
          default_zero(\$v3292\); default_zero(\$913\); 
          default_zero(\$1666_i\); default_zero(\$v1925\); 
          default_zero(\$v2310\); default_zero(\$v4012\); 
          default_zero(\$1616_lock\); default_zero(\$v2515\); 
          default_zero(\$v3545\); default_zero(\$v4175\); 
          default_zero(\$v3353\); default_zero(\$589\); 
          default_zero(\$v2157\); default_zero(\$v1835\); 
          default_zero(\$v3397\); default_zero(\$v4080\); 
          default_zero(\$v1681\); default_zero(\$805\); 
          default_zero(\$v2908\); default_zero(st); default_zero(\$v4138\); 
          default_zero(\$859\); default_zero(\$410\); default_zero(\$v29\); 
          default_zero(\$v60\); default_zero(\$v2325\); default_zero(\$860\); 
          default_zero(\$v3263\); default_zero(\$819\); default_zero(\$626\); 
          default_zero(\$1538\); default_zero(\$v58_lock\); 
          default_zero(\$1328\); default_zero(\$v3817\); 
          default_zero(\$v2686\); default_zero(\$v1617\); 
          default_zero(\$v77\); default_zero(\$v1934\); 
          default_zero(\$v4056\); default_zero(\$v3143\); 
          default_zero(\$489\); default_zero(\$709\); default_zero(\$v3727\); 
          default_zero(\$1494\); default_zero(\$v1716\); 
          default_zero(\$887\); default_zero(\$v1725\); 
          default_zero(\$v4220\); default_zero(\$1296\); 
          default_zero(\$v2961\); default_zero(\$v2235\); 
          default_zero(\$v1757\); default_zero(\$v4007\); 
          default_zero(\$809\); default_zero(\$1288\); default_zero(\$446\); 
          default_zero(\$1218\); default_zero(\$734_i\); 
          default_zero(\$v2834\); default_zero(\$354\); 
          default_zero(\$1027\); default_zero(\$292_i\); 
          default_zero(\$v102\); default_zero(\$v2920\); 
          default_zero(\$v2573\); default_zero(\$v3519\); 
          default_zero(\$1632\); default_zero(\$v3173\); 
          default_zero(\$1496\); default_zero(\$778_lock\); 
          default_zero(\$1487\); default_zero(\$499_lock\); 
          default_zero(\$v2699\); default_zero(\$v2312\); 
          default_zero(\$888\); default_zero(\$183_i\); 
          default_zero(\$v1543\); default_zero(\$919\); 
          default_zero(\$v1602\); default_zero(\$v1551\); 
          default_zero(\$v1871\); default_zero(\$1280\); 
          default_zero(\$752\); default_zero(\$570\); default_zero(\$v1915\); 
          default_zero(\$v3473\); default_zero(\$1124\); 
          default_zero(\$v3934\); default_zero(\$1262_lock\); 
          default_zero(\$409\); default_zero(\$v2649\); 
          default_zero(\$1427_lock\); default_zero(\$763\); 
          default_zero(\$635_i\); default_zero(\$242_lock\); 
          default_zero(\$v2910\); default_zero(\$1480\); 
          default_zero(\$839_x\); default_zero(\$1395\); 
          default_zero(\$240\); default_zero(\$v4228\); 
          default_zero(\$v1975\); default_zero(\$641\); 
          default_zero(\$1520\); default_zero(\$v3332\); 
          default_zero(\$1564\); default_zero(\$1573\); 
          default_zero(\$v2524\); default_zero(\$1463\); 
          default_zero(\$1159_lock\); default_zero(\$v2542\); 
          default_zero(\$v2879\); default_zero(\$v3878\); 
          default_zero(\$764_lock\); default_zero(\$215_lock\); 
          default_zero(\$505_lock\); default_zero(\$219\); 
          default_zero(\$1315_lock\); default_zero(\$533_lock\); 
          default_zero(\$329\); default_zero(\$661_lock\); 
          default_zero(\$v2339\); default_zero(\$359\); 
          default_zero(\$70_y\); default_zero(\$v2227\); 
          default_zero(\$v1863\); default_zero(\$1391\); 
          default_zero(\$v1592\); default_zero(\$625\); 
          default_zero(\$v4152\); default_zero(\$v2080\); 
          default_zero(\$1067\); default_zero(\$508\); 
          default_zero(\$v1574\); default_zero(\$v3055\); 
          default_zero(\$1281_lock\); default_zero(\$1684\); 
          default_zero(\$v2095\); default_zero(\$804_lock\); 
          default_zero(\$v3674\); default_zero(\$1235_lock\); 
          default_zero(\$v2052\); default_zero(\$1543\); 
          default_zero(\$v3849\); default_zero(\$846_lock\); 
          default_zero(\$1394\); default_zero(\$680\); 
          default_zero(\$179_lock\); default_zero(\$v18\); 
          default_zero(\$v2097\); default_zero(\$v2222\); 
          default_zero(\$v97\); default_zero(\$193\); default_zero(\$v3502\); 
          default_zero(\$1302\); default_zero(\$825\); 
          default_zero(\$v2474\); default_zero(\$1153\); 
          default_zero(\$1236_lock\); default_zero(\$453_lock\); 
          default_zero(\$v2607\); default_zero(\$1412\); 
          default_zero(\$1135\); default_zero(\$1130_lock\); 
          default_zero(\$v2730\); default_zero(\$411\); 
          default_zero(\$1509\); default_zero(\$v1672\); 
          default_zero(\$286\); default_zero(\$1396_x\); 
          default_zero(\$v3287\); default_zero(\$v2660\); 
          default_zero(\$v2210\); default_zero(\$1544\); 
          default_zero(\$v2075\); default_zero(\$178\); 
          default_zero(\$v1938\); default_zero(\$344\); 
          default_zero(\$v2482\); default_zero(\$1413\); 
          default_zero(\$1010_lock\); default_zero(\$v3019\); 
          default_zero(\$v2731\); default_zero(\$1538_lock\); 
          default_zero(\$345\); default_zero(\$1347\); default_zero(\$1160\); 
          default_zero(\$1371\); default_zero(\$v2617\); 
          default_zero(\$804\); default_zero(\$192_lock\); 
          default_zero(\$1166_lock\); default_zero(\$1355\); 
          default_zero(\$887_lock\); default_zero(\$v1611\); 
          default_zero(\$1620_i\); default_zero(\$617\); 
          default_zero(\$v2379\); default_zero(\$v1556\); 
          default_zero(\$v1836\); default_zero(\$v1916\); 
          default_zero(\$v1698\); default_zero(\$1615\); 
          default_zero(\$v39_lock\); default_zero(\$1353\); 
          default_zero(\$867_lock\); default_zero(\$v3432\); 
          default_zero(\$v98\); default_zero(\$814\); default_zero(\$v2501\); 
          rdy <= "1";
          rdy1455 := "0";
          \state\ <= compute1456;
          
        else if run = '1' then
          case \state\ is
          when \$147_forever1811388\ =>
            \state\ <= \$147_forever1811388\;
          when \$147_forever1811389\ =>
            \state\ <= \$147_forever1811389\;
          when \$147_forever1811390\ =>
            \state\ <= \$147_forever1811390\;
          when \$147_forever1811391\ =>
            \state\ <= \$147_forever1811391\;
          when \$147_forever1811392\ =>
            \state\ <= \$147_forever1811392\;
          when \$147_forever1811393\ =>
            \state\ <= \$147_forever1811393\;
          when \$147_forever1811394\ =>
            \state\ <= \$147_forever1811394\;
          when \$147_forever1811395\ =>
            \state\ <= \$147_forever1811395\;
          when \$147_forever1811396\ =>
            \state\ <= \$147_forever1811396\;
          when \$147_forever1811397\ =>
            \state\ <= \$147_forever1811397\;
          when \$147_forever1811398\ =>
            \state\ <= \$147_forever1811398\;
          when \$147_forever1811399\ =>
            \state\ <= \$147_forever1811399\;
          when \$147_forever1811400\ =>
            \state\ <= \$147_forever1811400\;
          when \$147_forever1811401\ =>
            \state\ <= \$147_forever1811401\;
          when \$147_forever1811402\ =>
            \state\ <= \$147_forever1811402\;
          when \$147_forever1811403\ =>
            \state\ <= \$147_forever1811403\;
          when \$147_forever1811404\ =>
            \state\ <= \$147_forever1811404\;
          when \$147_forever1811405\ =>
            \state\ <= \$147_forever1811405\;
          when \$147_forever1811406\ =>
            \state\ <= \$147_forever1811406\;
          when \$147_forever1811407\ =>
            \state\ <= \$147_forever1811407\;
          when \$147_forever1811408\ =>
            \state\ <= \$147_forever1811408\;
          when \$147_forever1811409\ =>
            \state\ <= \$147_forever1811409\;
          when \$147_forever1811410\ =>
            \state\ <= \$147_forever1811410\;
          when \$147_forever1811411\ =>
            \state\ <= \$147_forever1811411\;
          when \$147_forever1811412\ =>
            \state\ <= \$147_forever1811412\;
          when \$147_forever1811413\ =>
            \state\ <= \$147_forever1811413\;
          when \$147_forever1811414\ =>
            \state\ <= \$147_forever1811414\;
          when \$147_forever1811415\ =>
            \state\ <= \$147_forever1811415\;
          when \$147_forever1811416\ =>
            \state\ <= \$147_forever1811416\;
          when \$147_forever1811417\ =>
            \state\ <= \$147_forever1811417\;
          when \$147_forever1811418\ =>
            \state\ <= \$147_forever1811418\;
          when \$147_forever1811419\ =>
            \state\ <= \$147_forever1811419\;
          when \$147_forever1811420\ =>
            \state\ <= \$147_forever1811420\;
          when \$147_forever1811421\ =>
            \state\ <= \$147_forever1811421\;
          when \$147_forever1811422\ =>
            \state\ <= \$147_forever1811422\;
          when \$147_forever1811423\ =>
            \state\ <= \$147_forever1811423\;
          when \$147_forever1811424\ =>
            \state\ <= \$147_forever1811424\;
          when \$147_forever1811425\ =>
            \state\ <= \$147_forever1811425\;
          when \$147_forever1811426\ =>
            \state\ <= \$147_forever1811426\;
          when \$147_forever1811427\ =>
            \state\ <= \$147_forever1811427\;
          when \$147_forever1811428\ =>
            \state\ <= \$147_forever1811428\;
          when \$147_forever1811429\ =>
            \state\ <= \$147_forever1811429\;
          when \$147_forever1811430\ =>
            \state\ <= \$147_forever1811430\;
          when \$147_forever1811431\ =>
            \state\ <= \$147_forever1811431\;
          when \$147_forever1811432\ =>
            \state\ <= \$147_forever1811432\;
          when \$147_forever1811433\ =>
            \state\ <= \$147_forever1811433\;
          when \$147_forever1811434\ =>
            \state\ <= \$147_forever1811434\;
          when \$147_forever1811435\ =>
            \state\ <= \$147_forever1811435\;
          when \$147_forever1811436\ =>
            \state\ <= \$147_forever1811436\;
          when \$147_forever1811437\ =>
            \state\ <= \$147_forever1811437\;
          when \$147_forever1811438\ =>
            \state\ <= \$147_forever1811438\;
          when \$147_forever1811439\ =>
            \state\ <= \$147_forever1811439\;
          when \$147_forever1811440\ =>
            \state\ <= \$147_forever1811440\;
          when \$147_forever1811441\ =>
            \state\ <= \$147_forever1811441\;
          when \$147_forever1811442\ =>
            \state\ <= \$147_forever1811442\;
          when \$147_forever1811443\ =>
            \state\ <= \$147_forever1811443\;
          when \$147_forever1811444\ =>
            \state\ <= \$147_forever1811444\;
          when \$147_forever1811445\ =>
            \state\ <= \$147_forever1811445\;
          when \$147_forever1811446\ =>
            \state\ <= \$147_forever1811446\;
          when \$147_forever1811447\ =>
            \state\ <= \$147_forever1811447\;
          when \$147_forever1811448\ =>
            \state\ <= \$147_forever1811448\;
          when \$147_forever1811449\ =>
            \state\ <= \$147_forever1811449\;
          when \$147_forever1811450\ =>
            \state\ <= \$147_forever1811450\;
          when get_pause1462 =>
            \$v76_lock\ := eclat_false;
            \$v120\ := eclat_unit;
            \$v1460\ := \$arr1453_ptr_take\;
            if \$v1460\(0) = '1' then
              \state\ <= q_wait1459;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 17;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v120\;
              \state\ <= pause_setI1457;
            end if;
          when get_pause1479 =>
            \$v67_lock\ := eclat_false;
            \$v120\ := eclat_unit;
            \$v1460\ := \$arr1453_ptr_take\;
            if \$v1460\(0) = '1' then
              \state\ <= q_wait1459;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 17;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v120\;
              \state\ <= pause_setI1457;
            end if;
          when get_pause1504 =>
            \$v43_lock\ := eclat_false;
            \$70_y\ := \$84_x\;
            \$v1501\ := \$70_y\;
            \$v1502\ := \$v1501\(0 to 3);
            \$v1496\ := \$v1501\(4 to 35);
            case \$v1502\ is
            when "0001" =>
              a := \$v1496\(0 to 31);
              \$v1499\ := \$69_x\;
              \$v1500\ := \$v1499\(0 to 3);
              \$v1497\ := \$v1499\(4 to 35);
              case \$v1500\ is
              when "0001" =>
                b := \$v1497\(0 to 31);
                \$v1498\ := eclat_div(a & b);
                \$71_result_after_f\ := "0001" & \$v1498\;
                \$v1495\ := \$arr1452_ptr_take\;
                if \$v1495\(0) = '1' then
                  \state\ <= q_wait1494;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1492;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("* quotient arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811390\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("* quotient arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811389\;
            end case;
          when get_pause1572 =>
            \$180_lock\ := eclat_false;
            \$69_x\ := \$161_x\;
            \$v1570\ := \$arr1452_ptr_take\;
            if \$v1570\(0) = '1' then
              \state\ <= q_wait1569;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1567;
            end if;
          when get_pause1644 =>
            \$215_lock\ := eclat_false;
            \$v117\ := eclat_unit;
            \$v1642\ := \$arr1453_ptr_take\;
            if \$v1642\(0) = '1' then
              \state\ <= q_wait1641;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 16;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v117\;
              \state\ <= pause_setI1639;
            end if;
          when get_pause1661 =>
            \$214_lock\ := eclat_false;
            \$v117\ := eclat_unit;
            \$v1642\ := \$arr1453_ptr_take\;
            if \$v1642\(0) = '1' then
              \state\ <= q_wait1641;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 16;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v117\;
              \state\ <= pause_setI1639;
            end if;
          when get_pause1686 =>
            \$243_lock\ := eclat_false;
            \$208_y\ := \$224_x\;
            \$v1683\ := \$208_y\;
            \$v1684\ := \$v1683\(0 to 3);
            \$v1678\ := \$v1683\(4 to 35);
            case \$v1684\ is
            when "0001" =>
              \$26_a\ := \$v1678\(0 to 31);
              \$v1681\ := \$207_x\;
              \$v1682\ := \$v1681\(0 to 3);
              \$v1679\ := \$v1681\(4 to 35);
              case \$v1682\ is
              when "0001" =>
                b := \$v1679\(0 to 31);
                \$v1680\ := eclat_mult(\$26_a\ & b);
                \$209_result_after_f\ := "0001" & \$v1680\;
                \$v1677\ := \$arr1452_ptr_take\;
                if \$v1677\(0) = '1' then
                  \state\ <= q_wait1676;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1674;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("* arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811395\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("* arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811394\;
            end case;
          when get_pause1754 =>
            \$289_lock\ := eclat_false;
            \$207_x\ := \$270_x\;
            \$v1752\ := \$arr1452_ptr_take\;
            if \$v1752\(0) = '1' then
              \state\ <= q_wait1751;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1749;
            end if;
          when get_pause1826 =>
            \$324_lock\ := eclat_false;
            \$v114\ := eclat_unit;
            \$v1824\ := \$arr1453_ptr_take\;
            if \$v1824\(0) = '1' then
              \state\ <= q_wait1823;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 15;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v114\;
              \state\ <= pause_setI1821;
            end if;
          when get_pause1843 =>
            \$323_lock\ := eclat_false;
            \$v114\ := eclat_unit;
            \$v1824\ := \$arr1453_ptr_take\;
            if \$v1824\(0) = '1' then
              \state\ <= q_wait1823;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 15;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v114\;
              \state\ <= pause_setI1821;
            end if;
          when get_pause1868 =>
            \$352_lock\ := eclat_false;
            \$317_y\ := \$333_x\;
            \$v1865\ := \$317_y\;
            \$v1866\ := \$v1865\(0 to 3);
            \$v1860\ := \$v1865\(4 to 35);
            case \$v1866\ is
            when "0001" =>
              \$29_a\ := \$v1860\(0 to 31);
              \$v1863\ := \$316_x\;
              \$v1864\ := \$v1863\(0 to 3);
              \$v1861\ := \$v1863\(4 to 35);
              case \$v1864\ is
              when "0001" =>
                b := \$v1861\(0 to 31);
                \$v1862\ := eclat_sub(\$29_a\ & b);
                \$318_result_after_f\ := "0001" & \$v1862\;
                \$v1859\ := \$arr1452_ptr_take\;
                if \$v1859\(0) = '1' then
                  \state\ <= q_wait1858;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1856;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("- arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811400\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("- arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811399\;
            end case;
          when get_pause1936 =>
            \$398_lock\ := eclat_false;
            \$316_x\ := \$379_x\;
            \$v1934\ := \$arr1452_ptr_take\;
            if \$v1934\(0) = '1' then
              \state\ <= q_wait1933;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1931;
            end if;
          when get_pause2008 =>
            \$433_lock\ := eclat_false;
            \$v111\ := eclat_unit;
            \$v2006\ := \$arr1453_ptr_take\;
            if \$v2006\(0) = '1' then
              \state\ <= q_wait2005;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 14;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v111\;
              \state\ <= pause_setI2003;
            end if;
          when get_pause2025 =>
            \$432_lock\ := eclat_false;
            \$v111\ := eclat_unit;
            \$v2006\ := \$arr1453_ptr_take\;
            if \$v2006\(0) = '1' then
              \state\ <= q_wait2005;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 14;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v111\;
              \state\ <= pause_setI2003;
            end if;
          when get_pause2050 =>
            \$461_lock\ := eclat_false;
            \$426_y\ := \$442_x\;
            \$v2047\ := \$426_y\;
            \$v2048\ := \$v2047\(0 to 3);
            \$v2042\ := \$v2047\(4 to 35);
            case \$v2048\ is
            when "0001" =>
              \$32_a\ := \$v2042\(0 to 31);
              \$v2045\ := \$425_x\;
              \$v2046\ := \$v2045\(0 to 3);
              \$v2043\ := \$v2045\(4 to 35);
              case \$v2046\ is
              when "0001" =>
                b := \$v2043\(0 to 31);
                \$v2044\ := eclat_add(\$32_a\ & b);
                \$427_result_after_f\ := "0001" & \$v2044\;
                \$v2041\ := \$arr1452_ptr_take\;
                if \$v2041\(0) = '1' then
                  \state\ <= q_wait2040;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2038;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("+ arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811405\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("+ arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811404\;
            end case;
          when get_pause2118 =>
            \$507_lock\ := eclat_false;
            \$425_x\ := \$488_x\;
            \$v2116\ := \$arr1452_ptr_take\;
            if \$v2116\(0) = '1' then
              \state\ <= q_wait2115;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2113;
            end if;
          when get_pause2190 =>
            \$v58_lock\ := eclat_false;
            \$v108\ := eclat_unit;
            \$v2188\ := \$arr1453_ptr_take\;
            if \$v2188\(0) = '1' then
              \state\ <= q_wait2187;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 13;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v108\;
              \state\ <= pause_setI2185;
            end if;
          when get_pause2206 =>
            \$v55_lock\ := eclat_false;
            \$v108\ := eclat_unit;
            \$v2188\ := \$arr1453_ptr_take\;
            if \$v2188\(0) = '1' then
              \state\ <= q_wait2187;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 13;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v108\;
              \state\ <= pause_setI2185;
            end if;
          when get_pause2241 =>
            \$559_lock\ := eclat_false;
            \$53_y\ := \$540_x\;
            \$v2238\ := \$53_y\;
            \$v2239\ := \$v2238\(0 to 3);
            \$v2234\ := \$v2238\(4 to 35);
            case \$v2239\ is
            when "0001" =>
              \$35_a\ := \$v2234\(0 to 31);
              \$v2236\ := \$52_x\;
              \$v2237\ := \$v2236\(0 to 3);
              \$v2235\ := \$v2236\(4 to 35);
              case \$v2237\ is
              when "0001" =>
                b := \$v2235\(0 to 31);
                result := eclat_lt(\$35_a\ & b);
                \$v2233\ := \$arr1452_ptr_take\;
                if \$v2233\(0) = '1' then
                  \state\ <= q_wait2232;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2230;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("< arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811410\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("< arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811409\;
            end case;
          when get_pause2309 =>
            \$605_lock\ := eclat_false;
            \$52_x\ := \$586_x\;
            \$v2307\ := \$arr1452_ptr_take\;
            if \$v2307\(0) = '1' then
              \state\ <= q_wait2306;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2304;
            end if;
          when get_pause2381 =>
            \$640_lock\ := eclat_false;
            \$v106\ := eclat_unit;
            \$v2379\ := \$arr1453_ptr_take\;
            if \$v2379\(0) = '1' then
              \state\ <= q_wait2378;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 12;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v106\;
              \state\ <= pause_setI2376;
            end if;
          when get_pause2397 =>
            \$639_lock\ := eclat_false;
            \$v106\ := eclat_unit;
            \$v2379\ := \$arr1453_ptr_take\;
            if \$v2379\(0) = '1' then
              \state\ <= q_wait2378;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 12;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v106\;
              \state\ <= pause_setI2376;
            end if;
          when get_pause2435 =>
            \$661_lock\ := eclat_false;
            \$633_y\ := \$642_x\;
            \$v2432\ := \$633_y\;
            \$v2433\ := \$v2432\(0 to 3);
            \$v2425\ := \$v2432\(4 to 35);
            case \$v2433\ is
            when "0010" =>
              ta := \$v2425\(0 to 31);
              \$v2427\ := \$632_x\;
              \$v2428\ := \$v2427\(0 to 3);
              \$v2426\ := \$v2427\(4 to 35);
              case \$v2428\ is
              when "0010" =>
                tb := \$v2426\(0 to 31);
                \$634_result\ := eclat_eq(ta & tb);
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              when others =>
                \$634_result\ := eclat_false;
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              end case;
            when "0001" =>
              ia := \$v2425\(0 to 31);
              \$v2430\ := \$632_x\;
              \$v2431\ := \$v2430\(0 to 3);
              \$v2429\ := \$v2430\(4 to 35);
              case \$v2431\ is
              when "0001" =>
                ib := \$v2429\(0 to 31);
                \$634_result\ := eclat_eq(ia & ib);
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              when others =>
                \$634_result\ := eclat_false;
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              end case;
            when others =>
              \$634_result\ := eclat_false;
              \$v2424\ := \$arr1452_ptr_take\;
              if \$v2424\(0) = '1' then
                \state\ <= q_wait2423;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2421;
              end if;
            end case;
          when get_pause2503 =>
            \$707_lock\ := eclat_false;
            \$632_x\ := \$688_x\;
            \$v2501\ := \$arr1452_ptr_take\;
            if \$v2501\(0) = '1' then
              \state\ <= q_wait2500;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2498;
            end if;
          when get_pause2575 =>
            \$739_lock\ := eclat_false;
            \$v104\ := eclat_unit;
            \$v2573\ := \$arr1453_ptr_take\;
            if \$v2573\(0) = '1' then
              \state\ <= q_wait2572;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 11;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v104\;
              \state\ <= pause_setI2570;
            end if;
          when get_pause2585 =>
            \$738_lock\ := eclat_false;
            \$v104\ := eclat_unit;
            \$v2573\ := \$arr1453_ptr_take\;
            if \$v2573\(0) = '1' then
              \state\ <= q_wait2572;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 11;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v104\;
              \state\ <= pause_setI2570;
            end if;
          when get_pause2615 =>
            \$766_lock\ := eclat_false;
            \$83_x\ := \$747_x\;
            \$v2612\ := \$83_x\;
            \$v2613\ := \$v2612\(0 to 3);
            \$v2607\ := \$v2612\(4 to 35);
            case \$v2613\ is
            when "0010" =>
              \$135_i\ := \$v2607\(0 to 31);
              \$v2611\ := \$arr1451_ptr_take\;
              if \$v2611\(0) = '1' then
                \state\ <= q_wait2610;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$135_i\));
                \state\ <= pause_getI2608;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811417\;
            end case;
          when get_pause2683 =>
            \$812_lock\ := eclat_false;
            \$55_x\ := \$793_x\;
            \$v2681\ := \$arr1452_ptr_take\;
            if \$v2681\(0) = '1' then
              \state\ <= q_wait2680;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2678;
            end if;
          when get_pause2755 =>
            \$846_lock\ := eclat_false;
            \$v102\ := eclat_unit;
            \$v2753\ := \$arr1453_ptr_take\;
            if \$v2753\(0) = '1' then
              \state\ <= q_wait2752;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 10;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v102\;
              \state\ <= pause_setI2750;
            end if;
          when get_pause2765 =>
            \$845_lock\ := eclat_false;
            \$v102\ := eclat_unit;
            \$v2753\ := \$arr1453_ptr_take\;
            if \$v2753\(0) = '1' then
              \state\ <= q_wait2752;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 10;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v102\;
              \state\ <= pause_setI2750;
            end if;
          when get_pause2795 =>
            \$875_lock\ := eclat_false;
            \$851_x\ := \$856_x\;
            \$v2792\ := \$851_x\;
            \$v2793\ := \$v2792\(0 to 3);
            \$v2787\ := \$v2792\(4 to 35);
            case \$v2793\ is
            when "0010" =>
              \$852_i\ := \$v2787\(0 to 31);
              \$v2791\ := \$arr1451_ptr_take\;
              if \$v2791\(0) = '1' then
                \state\ <= q_wait2790;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$852_i\));
                \state\ <= pause_getI2788;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811421\;
            end case;
          when get_pause2863 =>
            \$921_lock\ := eclat_false;
            \$839_x\ := \$902_x\;
            \$v2861\ := \$arr1452_ptr_take\;
            if \$v2861\(0) = '1' then
              \state\ <= q_wait2860;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2858;
            end if;
          when get_pause2935 =>
            \$955_lock\ := eclat_false;
            \$v100\ := eclat_unit;
            \$v2933\ := \$arr1453_ptr_take\;
            if \$v2933\(0) = '1' then
              \state\ <= q_wait2932;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 9;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v100\;
              \state\ <= pause_setI2930;
            end if;
          when get_pause2945 =>
            \$954_lock\ := eclat_false;
            \$v100\ := eclat_unit;
            \$v2933\ := \$arr1453_ptr_take\;
            if \$v2933\(0) = '1' then
              \state\ <= q_wait2932;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 9;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v100\;
              \state\ <= pause_setI2930;
            end if;
          when get_pause2975 =>
            \$984_lock\ := eclat_false;
            \$960_x\ := \$965_x\;
            \$v2972\ := \$960_x\;
            \$v2973\ := \$v2972\(0 to 3);
            \$v2967\ := \$v2972\(4 to 35);
            case \$v2973\ is
            when "0010" =>
              \$961_i\ := \$v2967\(0 to 31);
              \$v2971\ := \$arr1451_ptr_take\;
              if \$v2971\(0) = '1' then
                \state\ <= q_wait2970;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$961_i\));
                \state\ <= pause_getI2968;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811425\;
            end case;
          when get_pause3043 =>
            \$1030_lock\ := eclat_false;
            \$948_x\ := \$1011_x\;
            \$v3041\ := \$arr1452_ptr_take\;
            if \$v3041\(0) = '1' then
              \state\ <= q_wait3040;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3038;
            end if;
          when get_pause3115 =>
            \$1065_lock\ := eclat_false;
            \$v98\ := eclat_unit;
            \$v3113\ := \$arr1453_ptr_take\;
            if \$v3113\(0) = '1' then
              \state\ <= q_wait3112;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 8;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v98\;
              \state\ <= pause_setI3110;
            end if;
          when get_pause3132 =>
            \$1061_lock\ := eclat_false;
            \$v98\ := eclat_unit;
            \$v3113\ := \$arr1453_ptr_take\;
            if \$v3113\(0) = '1' then
              \state\ <= q_wait3112;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 8;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v98\;
              \state\ <= pause_setI3110;
            end if;
          when get_pause3157 =>
            \$1098_lock\ := eclat_false;
            \$1074_x\ := \$1079_x\;
            \$v3154\ := \$1074_x\;
            \$v3155\ := \$v3154\(0 to 3);
            \$v3149\ := \$v3154\(4 to 35);
            case \$v3155\ is
            when "0010" =>
              \$1075_i\ := \$v3149\(0 to 31);
              \$v3153\ := \$arr1451_ptr_take\;
              if \$v3153\(0) = '1' then
                \state\ <= q_wait3152;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1075_i\));
                \state\ <= pause_getI3150;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811429\;
            end case;
          when get_pause3229 =>
            \$1134_lock\ := eclat_false;
            \$v97\ := eclat_unit;
            \$v3227\ := \$arr1453_ptr_take\;
            if \$v3227\(0) = '1' then
              \state\ <= q_wait3226;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 7;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v97\;
              \state\ <= pause_setI3224;
            end if;
          when get_pause3246 =>
            \$1130_lock\ := eclat_false;
            \$v97\ := eclat_unit;
            \$v3227\ := \$arr1453_ptr_take\;
            if \$v3227\(0) = '1' then
              \state\ <= q_wait3226;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 7;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v97\;
              \state\ <= pause_setI3224;
            end if;
          when get_pause3271 =>
            \$1167_lock\ := eclat_false;
            \$1143_x\ := \$1148_x\;
            \$v3268\ := \$1143_x\;
            \$v3269\ := \$v3268\(0 to 3);
            \$v3263\ := \$v3268\(4 to 35);
            case \$v3269\ is
            when "0010" =>
              \$1144_i\ := \$v3263\(0 to 31);
              \$v3267\ := \$arr1451_ptr_take\;
              if \$v3267\(0) = '1' then
                \state\ <= q_wait3266;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1144_i\));
                \state\ <= pause_getI3264;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811432\;
            end case;
          when get_pause3343 =>
            \$1203_lock\ := eclat_false;
            \$v96\ := eclat_unit;
            \$v3341\ := \$arr1453_ptr_take\;
            if \$v3341\(0) = '1' then
              \state\ <= q_wait3340;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 6;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v96\;
              \state\ <= pause_setI3338;
            end if;
          when get_pause3360 =>
            \$1199_lock\ := eclat_false;
            \$v96\ := eclat_unit;
            \$v3341\ := \$arr1453_ptr_take\;
            if \$v3341\(0) = '1' then
              \state\ <= q_wait3340;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 6;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v96\;
              \state\ <= pause_setI3338;
            end if;
          when get_pause3385 =>
            \$1236_lock\ := eclat_false;
            \$1212_x\ := \$1217_x\;
            \$v3382\ := \$1212_x\;
            \$v3383\ := \$v3382\(0 to 3);
            \$v3377\ := \$v3382\(4 to 35);
            case \$v3383\ is
            when "0010" =>
              \$1213_i\ := \$v3377\(0 to 31);
              \$v3381\ := \$arr1451_ptr_take\;
              if \$v3381\(0) = '1' then
                \state\ <= q_wait3380;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1213_i\));
                \state\ <= pause_getI3378;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811435\;
            end case;
          when get_pause3457 =>
            \$1268_lock\ := eclat_false;
            \$v95\ := eclat_unit;
            \$v3455\ := \$arr1453_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 5;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v95\;
              \state\ <= pause_setI3452;
            end if;
          when get_pause3467 =>
            \$1267_lock\ := eclat_false;
            \$v95\ := eclat_unit;
            \$v3455\ := \$arr1453_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 5;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v95\;
              \state\ <= pause_setI3452;
            end if;
          when get_pause3499 =>
            \$1289_lock\ := eclat_false;
            \$73_result\ := \$1270_x\;
            \$v3496\ := \$73_result\;
            \$v3497\ := \$v3496\(0 to 3);
            \$v3489\ := \$v3496\(4 to 35);
            case \$v3497\ is
            when "0010" =>
              \$v3490\ := "00000000000000000000000000000000";
              \$v3491\ := "00000000000000000000000000000000";
              \$v3492\ := "00000000000000000000000000000101";
              \$74_result_after_f\ := "0001" & \$v3490\ & "0001" & \$v3491\ & "0001" & \$v3492\;
              \$v3488\ := \$arr1452_ptr_take\;
              if \$v3488\(0) = '1' then
                \state\ <= q_wait3487;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3485;
              end if;
            when others =>
              \$v3493\ := "00000000000000000000000000000001";
              \$v3494\ := "00000000000000000000000000000010";
              \$v3495\ := "00000000000000000000000000000101";
              \$74_result_after_f\ := "0010" & \$v3493\ & "0010" & \$v3494\ & "0001" & \$v3495\;
              \$v3488\ := \$arr1452_ptr_take\;
              if \$v3488\(0) = '1' then
                \state\ <= q_wait3487;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3485;
              end if;
            end case;
          when get_pause3571 =>
            \$1324_lock\ := eclat_false;
            \$v94\ := eclat_unit;
            \$v3569\ := \$arr1453_ptr_take\;
            if \$v3569\(0) = '1' then
              \state\ <= q_wait3568;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 4;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v94\;
              \state\ <= pause_setI3566;
            end if;
          when get_pause3582 =>
            \$1320_lock\ := eclat_false;
            \$v94\ := eclat_unit;
            \$v3569\ := \$arr1453_ptr_take\;
            if \$v3569\(0) = '1' then
              \state\ <= q_wait3568;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 4;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v94\;
              \state\ <= pause_setI3566;
            end if;
          when get_pause3622 =>
            \$1356_lock\ := eclat_false;
            \$1332_x\ := \$1337_x\;
            \$v3619\ := \$1332_x\;
            \$v3620\ := \$v3619\(0 to 3);
            \$v3614\ := \$v3619\(4 to 35);
            case \$v3620\ is
            when "0010" =>
              \$1333_i\ := \$v3614\(0 to 31);
              \$v3618\ := \$arr1451_ptr_take\;
              if \$v3618\(0) = '1' then
                \state\ <= q_wait3617;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1333_i\));
                \state\ <= pause_getI3615;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811440\;
            end case;
          when get_pause3694 =>
            \$1390_lock\ := eclat_false;
            \$v93\ := eclat_unit;
            \$v3692\ := \$arr1453_ptr_take\;
            if \$v3692\(0) = '1' then
              \state\ <= q_wait3691;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 3;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v93\;
              \state\ <= pause_setI3689;
            end if;
          when get_pause3711 =>
            \$1389_lock\ := eclat_false;
            \$v93\ := eclat_unit;
            \$v3692\ := \$arr1453_ptr_take\;
            if \$v3692\(0) = '1' then
              \state\ <= q_wait3691;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 3;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v93\;
              \state\ <= pause_setI3689;
            end if;
          when get_pause3729 =>
            \$1415_lock\ := eclat_false;
            \$v3727\ := \$arr1452_ptr_take\;
            if \$v3727\(0) = '1' then
              \state\ <= q_wait3726;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3724;
            end if;
          when get_pause3797 =>
            \$1461_lock\ := eclat_false;
            \$1383_x\ := \$1442_x\;
            \$v3795\ := \$arr1452_ptr_take\;
            if \$v3795\(0) = '1' then
              \state\ <= q_wait3794;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3792;
            end if;
          when get_pause3869 =>
            \$1493_lock\ := eclat_false;
            \$v91\ := eclat_unit;
            \$v3867\ := \$arr1453_ptr_take\;
            if \$v3867\(0) = '1' then
              \state\ <= q_wait3866;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 1;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v91\;
              \state\ <= pause_setI3864;
            end if;
          when get_pause3886 =>
            \$1492_lock\ := eclat_false;
            \$v91\ := eclat_unit;
            \$v3867\ := \$arr1453_ptr_take\;
            if \$v3867\(0) = '1' then
              \state\ <= q_wait3866;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 1;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v91\;
              \state\ <= pause_setI3864;
            end if;
          when get_pause3904 =>
            \$1518_lock\ := eclat_false;
            \$76_result\ := \$1499_x\;
            \$v3902\ := \$arr1452_ptr_take\;
            if \$v3902\(0) = '1' then
              \state\ <= q_wait3901;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3899;
            end if;
          when get_pause3976 =>
            \$1550_lock\ := eclat_false;
            \$v89\ := eclat_unit;
            \$v3974\ := \$arr1453_ptr_take\;
            if \$v3974\(0) = '1' then
              \state\ <= q_wait3973;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 0;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v89\;
              \state\ <= pause_setI3971;
            end if;
          when get_pause3986 =>
            \$1549_lock\ := eclat_false;
            \$v89\ := eclat_unit;
            \$v3974\ := \$arr1453_ptr_take\;
            if \$v3974\(0) = '1' then
              \state\ <= q_wait3973;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 0;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v89\;
              \state\ <= pause_setI3971;
            end if;
          when get_pause4009 =>
            \$1571_lock\ := eclat_false;
            \$67_z\ := \$1552_x\;
            \$v4007\ := \$arr1452_ptr_take\;
            if \$v4007\(0) = '1' then
              \state\ <= q_wait4006;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4004;
            end if;
          when get_pause4077 =>
            \$1617_lock\ := eclat_false;
            \$66_y\ := \$1598_x\;
            \$v4075\ := \$arr1452_ptr_take\;
            if \$v4075\(0) = '1' then
              \state\ <= q_wait4074;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4072;
            end if;
          when get_pause4145 =>
            \$1663_lock\ := eclat_false;
            \$65_x\ := \$1644_x\;
            \$v4143\ := \$arr1452_ptr_take\;
            if \$v4143\(0) = '1' then
              \state\ <= q_wait4142;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4140;
            end if;
          when get_wait1461 =>
            if \$v76_lock\(0) = '1' then
              \state\ <= get_wait1461;
            else
              \$v76_lock\ := eclat_true;
              \state\ <= get_pause1462;
            end if;
          when get_wait1463 =>
            if \$v73_lock\(0) = '1' then
              \state\ <= get_wait1463;
            else
              \$v74\ := \$v73\;
              \$v75\ := \$v74\ & "00000000000000000000000000000001";
              \$v77\ := eclat_sub(\$v75\);
              if \$v76_lock\(0) = '1' then
                \state\ <= get_wait1461;
              else
                \$v76_lock\ := eclat_true;
                \state\ <= get_pause1462;
              end if;
            end if;
          when get_wait1478 =>
            if \$v67_lock\(0) = '1' then
              \state\ <= get_wait1478;
            else
              \$v67_lock\ := eclat_true;
              \state\ <= get_pause1479;
            end if;
          when get_wait1491 =>
            if \$v60_lock\(0) = '1' then
              \state\ <= get_wait1491;
            else
              \$81_i\ := \$v60\;
              \$v1490\ := eclat_gt(\$81_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1490\(0) = '1' then
                \$v1489\ := eclat_eq(\$81_i\ & X"000" & X"15f90");
                if \$v1489\(0) = '1' then
                  \$v1477\ := \$arr1451_ptr_take\;
                  if \$v1477\(0) = '1' then
                    \state\ <= q_wait1476;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1472\ := "00000000000000000000000000000000";
                    \$v1473\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$71_result_after_f\ & "0001" & \$v1472\ & "0001" & \$v1473\;
                    \state\ <= pause_setI1474;
                  end if;
                else
                  \$v1488\ := \$arr1451_ptr_take\;
                  if \$v1488\(0) = '1' then
                    \state\ <= q_wait1487;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1484\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$71_result_after_f\ & "0010" & \$81_i\ & "0001" & \$v1484\;
                    \state\ <= pause_setI1485;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811388\;
              end if;
            end if;
          when get_wait1503 =>
            if \$v43_lock\(0) = '1' then
              \state\ <= get_wait1503;
            else
              \$v43_lock\ := eclat_true;
              \state\ <= get_pause1504;
            end if;
          when get_wait1512 =>
            if \$v39_lock\(0) = '1' then
              \state\ <= get_wait1512;
            else
              \$v40\ := \$v39\;
              \$v1511\ := \$arr1451_ptr_take\;
              if \$v1511\(0) = '1' then
                \state\ <= q_wait1510;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v40\));
                \state\ <= pause_getI1508;
              end if;
            end if;
          when get_wait1530 =>
            if \$v31_lock\(0) = '1' then
              \state\ <= get_wait1530;
            else
              \$v32\ := \$v31\;
              \$v1529\ := \$arr1451_ptr_take\;
              if \$v1529\(0) = '1' then
                \state\ <= q_wait1528;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v32\));
                \state\ <= pause_getI1526;
              end if;
            end if;
          when get_wait1539 =>
            if \$v28_lock\(0) = '1' then
              \state\ <= get_wait1539;
            else
              \$v29\ := \$v28\;
              \$v1538\ := \$arr1451_ptr_take\;
              if \$v1538\(0) = '1' then
                \state\ <= q_wait1537;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v29\));
                \state\ <= pause_getI1535;
              end if;
            end if;
          when get_wait1544 =>
            if \$v27_lock\(0) = '1' then
              \state\ <= get_wait1544;
            else
              \$v37\ := \$v27\;
              \$v1543\ := \$arr1452_ptr_take\;
              if \$v1543\(0) = '1' then
                \state\ <= q_wait1542;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1540;
              end if;
            end if;
          when get_wait1557 =>
            if \$v22_lock\(0) = '1' then
              \state\ <= get_wait1557;
            else
              \$v23\ := \$v22\;
              \$v1556\ := \$arr1451_ptr_take\;
              if \$v1556\(0) = '1' then
                \state\ <= q_wait1555;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v23\));
                \state\ <= pause_getI1553;
              end if;
            end if;
          when get_wait1566 =>
            if \$v19_lock\(0) = '1' then
              \state\ <= get_wait1566;
            else
              \$v20\ := \$v19\;
              \$v1565\ := \$arr1451_ptr_take\;
              if \$v1565\(0) = '1' then
                \state\ <= q_wait1564;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v20\));
                \state\ <= pause_getI1562;
              end if;
            end if;
          when get_wait1571 =>
            if \$180_lock\(0) = '1' then
              \state\ <= get_wait1571;
            else
              \$180_lock\ := eclat_true;
              \state\ <= get_pause1572;
            end if;
          when get_wait1580 =>
            if \$192_lock\(0) = '1' then
              \state\ <= get_wait1580;
            else
              \$191\ := \$192\;
              \$v1579\ := \$arr1451_ptr_take\;
              if \$v1579\(0) = '1' then
                \state\ <= q_wait1578;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$191\));
                \state\ <= pause_getI1576;
              end if;
            end if;
          when get_wait1598 =>
            if \$172_lock\(0) = '1' then
              \state\ <= get_wait1598;
            else
              \$171\ := \$172\;
              \$v1597\ := \$arr1451_ptr_take\;
              if \$v1597\(0) = '1' then
                \state\ <= q_wait1596;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$171\));
                \state\ <= pause_getI1594;
              end if;
            end if;
          when get_wait1607 =>
            if \$178_lock\(0) = '1' then
              \state\ <= get_wait1607;
            else
              \$177\ := \$178\;
              \$v1606\ := \$arr1451_ptr_take\;
              if \$v1606\(0) = '1' then
                \state\ <= q_wait1605;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$177\));
                \state\ <= pause_getI1603;
              end if;
            end if;
          when get_wait1612 =>
            if \$179_lock\(0) = '1' then
              \state\ <= get_wait1612;
            else
              \$163\ := \$179\;
              \$v1611\ := \$arr1452_ptr_take\;
              if \$v1611\(0) = '1' then
                \state\ <= q_wait1610;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1608;
              end if;
            end if;
          when get_wait1625 =>
            if \$200_lock\(0) = '1' then
              \state\ <= get_wait1625;
            else
              \$199\ := \$200\;
              \$v1624\ := \$arr1451_ptr_take\;
              if \$v1624\(0) = '1' then
                \state\ <= q_wait1623;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$199\));
                \state\ <= pause_getI1621;
              end if;
            end if;
          when get_wait1634 =>
            if \$206_lock\(0) = '1' then
              \state\ <= get_wait1634;
            else
              \$205\ := \$206\;
              \$v1633\ := \$arr1451_ptr_take\;
              if \$v1633\(0) = '1' then
                \state\ <= q_wait1632;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$205\));
                \state\ <= pause_getI1630;
              end if;
            end if;
          when get_wait1643 =>
            if \$215_lock\(0) = '1' then
              \state\ <= get_wait1643;
            else
              \$215_lock\ := eclat_true;
              \state\ <= get_pause1644;
            end if;
          when get_wait1645 =>
            if \$219_lock\(0) = '1' then
              \state\ <= get_wait1645;
            else
              \$218\ := \$219\;
              \$217\ := \$218\ & "00000000000000000000000000000001";
              \$216\ := eclat_sub(\$217\);
              if \$215_lock\(0) = '1' then
                \state\ <= get_wait1643;
              else
                \$215_lock\ := eclat_true;
                \state\ <= get_pause1644;
              end if;
            end if;
          when get_wait1660 =>
            if \$214_lock\(0) = '1' then
              \state\ <= get_wait1660;
            else
              \$214_lock\ := eclat_true;
              \state\ <= get_pause1661;
            end if;
          when get_wait1673 =>
            if \$220_lock\(0) = '1' then
              \state\ <= get_wait1673;
            else
              \$210_i\ := \$220\;
              \$v1672\ := eclat_gt(\$210_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1672\(0) = '1' then
                \$v1671\ := eclat_eq(\$210_i\ & X"000" & X"15f90");
                if \$v1671\(0) = '1' then
                  \$v1659\ := \$arr1451_ptr_take\;
                  if \$v1659\(0) = '1' then
                    \state\ <= q_wait1658;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1654\ := "00000000000000000000000000000000";
                    \$v1655\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$209_result_after_f\ & "0001" & \$v1654\ & "0001" & \$v1655\;
                    \state\ <= pause_setI1656;
                  end if;
                else
                  \$v1670\ := \$arr1451_ptr_take\;
                  if \$v1670\(0) = '1' then
                    \state\ <= q_wait1669;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1666\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$209_result_after_f\ & "0010" & \$210_i\ & "0001" & \$v1666\;
                    \state\ <= pause_setI1667;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811393\;
              end if;
            end if;
          when get_wait1685 =>
            if \$243_lock\(0) = '1' then
              \state\ <= get_wait1685;
            else
              \$243_lock\ := eclat_true;
              \state\ <= get_pause1686;
            end if;
          when get_wait1694 =>
            if \$255_lock\(0) = '1' then
              \state\ <= get_wait1694;
            else
              \$254\ := \$255\;
              \$v1693\ := \$arr1451_ptr_take\;
              if \$v1693\(0) = '1' then
                \state\ <= q_wait1692;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$254\));
                \state\ <= pause_getI1690;
              end if;
            end if;
          when get_wait1712 =>
            if \$235_lock\(0) = '1' then
              \state\ <= get_wait1712;
            else
              \$234\ := \$235\;
              \$v1711\ := \$arr1451_ptr_take\;
              if \$v1711\(0) = '1' then
                \state\ <= q_wait1710;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$234\));
                \state\ <= pause_getI1708;
              end if;
            end if;
          when get_wait1721 =>
            if \$241_lock\(0) = '1' then
              \state\ <= get_wait1721;
            else
              \$240\ := \$241\;
              \$v1720\ := \$arr1451_ptr_take\;
              if \$v1720\(0) = '1' then
                \state\ <= q_wait1719;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$240\));
                \state\ <= pause_getI1717;
              end if;
            end if;
          when get_wait1726 =>
            if \$242_lock\(0) = '1' then
              \state\ <= get_wait1726;
            else
              \$226\ := \$242\;
              \$v1725\ := \$arr1452_ptr_take\;
              if \$v1725\(0) = '1' then
                \state\ <= q_wait1724;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1722;
              end if;
            end if;
          when get_wait1739 =>
            if \$263_lock\(0) = '1' then
              \state\ <= get_wait1739;
            else
              \$262\ := \$263\;
              \$v1738\ := \$arr1451_ptr_take\;
              if \$v1738\(0) = '1' then
                \state\ <= q_wait1737;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$262\));
                \state\ <= pause_getI1735;
              end if;
            end if;
          when get_wait1748 =>
            if \$269_lock\(0) = '1' then
              \state\ <= get_wait1748;
            else
              \$268\ := \$269\;
              \$v1747\ := \$arr1451_ptr_take\;
              if \$v1747\(0) = '1' then
                \state\ <= q_wait1746;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$268\));
                \state\ <= pause_getI1744;
              end if;
            end if;
          when get_wait1753 =>
            if \$289_lock\(0) = '1' then
              \state\ <= get_wait1753;
            else
              \$289_lock\ := eclat_true;
              \state\ <= get_pause1754;
            end if;
          when get_wait1762 =>
            if \$301_lock\(0) = '1' then
              \state\ <= get_wait1762;
            else
              \$300\ := \$301\;
              \$v1761\ := \$arr1451_ptr_take\;
              if \$v1761\(0) = '1' then
                \state\ <= q_wait1760;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$300\));
                \state\ <= pause_getI1758;
              end if;
            end if;
          when get_wait1780 =>
            if \$281_lock\(0) = '1' then
              \state\ <= get_wait1780;
            else
              \$280\ := \$281\;
              \$v1779\ := \$arr1451_ptr_take\;
              if \$v1779\(0) = '1' then
                \state\ <= q_wait1778;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$280\));
                \state\ <= pause_getI1776;
              end if;
            end if;
          when get_wait1789 =>
            if \$287_lock\(0) = '1' then
              \state\ <= get_wait1789;
            else
              \$286\ := \$287\;
              \$v1788\ := \$arr1451_ptr_take\;
              if \$v1788\(0) = '1' then
                \state\ <= q_wait1787;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$286\));
                \state\ <= pause_getI1785;
              end if;
            end if;
          when get_wait1794 =>
            if \$288_lock\(0) = '1' then
              \state\ <= get_wait1794;
            else
              \$272\ := \$288\;
              \$v1793\ := \$arr1452_ptr_take\;
              if \$v1793\(0) = '1' then
                \state\ <= q_wait1792;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1790;
              end if;
            end if;
          when get_wait1807 =>
            if \$309_lock\(0) = '1' then
              \state\ <= get_wait1807;
            else
              \$308\ := \$309\;
              \$v1806\ := \$arr1451_ptr_take\;
              if \$v1806\(0) = '1' then
                \state\ <= q_wait1805;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$308\));
                \state\ <= pause_getI1803;
              end if;
            end if;
          when get_wait1816 =>
            if \$315_lock\(0) = '1' then
              \state\ <= get_wait1816;
            else
              \$314\ := \$315\;
              \$v1815\ := \$arr1451_ptr_take\;
              if \$v1815\(0) = '1' then
                \state\ <= q_wait1814;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$314\));
                \state\ <= pause_getI1812;
              end if;
            end if;
          when get_wait1825 =>
            if \$324_lock\(0) = '1' then
              \state\ <= get_wait1825;
            else
              \$324_lock\ := eclat_true;
              \state\ <= get_pause1826;
            end if;
          when get_wait1827 =>
            if \$328_lock\(0) = '1' then
              \state\ <= get_wait1827;
            else
              \$327\ := \$328\;
              \$326\ := \$327\ & "00000000000000000000000000000001";
              \$325\ := eclat_sub(\$326\);
              if \$324_lock\(0) = '1' then
                \state\ <= get_wait1825;
              else
                \$324_lock\ := eclat_true;
                \state\ <= get_pause1826;
              end if;
            end if;
          when get_wait1842 =>
            if \$323_lock\(0) = '1' then
              \state\ <= get_wait1842;
            else
              \$323_lock\ := eclat_true;
              \state\ <= get_pause1843;
            end if;
          when get_wait1855 =>
            if \$329_lock\(0) = '1' then
              \state\ <= get_wait1855;
            else
              \$319_i\ := \$329\;
              \$v1854\ := eclat_gt(\$319_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1854\(0) = '1' then
                \$v1853\ := eclat_eq(\$319_i\ & X"000" & X"15f90");
                if \$v1853\(0) = '1' then
                  \$v1841\ := \$arr1451_ptr_take\;
                  if \$v1841\(0) = '1' then
                    \state\ <= q_wait1840;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1836\ := "00000000000000000000000000000000";
                    \$v1837\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$318_result_after_f\ & "0001" & \$v1836\ & "0001" & \$v1837\;
                    \state\ <= pause_setI1838;
                  end if;
                else
                  \$v1852\ := \$arr1451_ptr_take\;
                  if \$v1852\(0) = '1' then
                    \state\ <= q_wait1851;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1848\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$318_result_after_f\ & "0010" & \$319_i\ & "0001" & \$v1848\;
                    \state\ <= pause_setI1849;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811398\;
              end if;
            end if;
          when get_wait1867 =>
            if \$352_lock\(0) = '1' then
              \state\ <= get_wait1867;
            else
              \$352_lock\ := eclat_true;
              \state\ <= get_pause1868;
            end if;
          when get_wait1876 =>
            if \$364_lock\(0) = '1' then
              \state\ <= get_wait1876;
            else
              \$363\ := \$364\;
              \$v1875\ := \$arr1451_ptr_take\;
              if \$v1875\(0) = '1' then
                \state\ <= q_wait1874;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$363\));
                \state\ <= pause_getI1872;
              end if;
            end if;
          when get_wait1894 =>
            if \$344_lock\(0) = '1' then
              \state\ <= get_wait1894;
            else
              \$343\ := \$344\;
              \$v1893\ := \$arr1451_ptr_take\;
              if \$v1893\(0) = '1' then
                \state\ <= q_wait1892;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$343\));
                \state\ <= pause_getI1890;
              end if;
            end if;
          when get_wait1903 =>
            if \$350_lock\(0) = '1' then
              \state\ <= get_wait1903;
            else
              \$349\ := \$350\;
              \$v1902\ := \$arr1451_ptr_take\;
              if \$v1902\(0) = '1' then
                \state\ <= q_wait1901;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$349\));
                \state\ <= pause_getI1899;
              end if;
            end if;
          when get_wait1908 =>
            if \$351_lock\(0) = '1' then
              \state\ <= get_wait1908;
            else
              \$335\ := \$351\;
              \$v1907\ := \$arr1452_ptr_take\;
              if \$v1907\(0) = '1' then
                \state\ <= q_wait1906;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1904;
              end if;
            end if;
          when get_wait1921 =>
            if \$372_lock\(0) = '1' then
              \state\ <= get_wait1921;
            else
              \$371\ := \$372\;
              \$v1920\ := \$arr1451_ptr_take\;
              if \$v1920\(0) = '1' then
                \state\ <= q_wait1919;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$371\));
                \state\ <= pause_getI1917;
              end if;
            end if;
          when get_wait1930 =>
            if \$378_lock\(0) = '1' then
              \state\ <= get_wait1930;
            else
              \$377\ := \$378\;
              \$v1929\ := \$arr1451_ptr_take\;
              if \$v1929\(0) = '1' then
                \state\ <= q_wait1928;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$377\));
                \state\ <= pause_getI1926;
              end if;
            end if;
          when get_wait1935 =>
            if \$398_lock\(0) = '1' then
              \state\ <= get_wait1935;
            else
              \$398_lock\ := eclat_true;
              \state\ <= get_pause1936;
            end if;
          when get_wait1944 =>
            if \$410_lock\(0) = '1' then
              \state\ <= get_wait1944;
            else
              \$409\ := \$410\;
              \$v1943\ := \$arr1451_ptr_take\;
              if \$v1943\(0) = '1' then
                \state\ <= q_wait1942;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$409\));
                \state\ <= pause_getI1940;
              end if;
            end if;
          when get_wait1962 =>
            if \$390_lock\(0) = '1' then
              \state\ <= get_wait1962;
            else
              \$389\ := \$390\;
              \$v1961\ := \$arr1451_ptr_take\;
              if \$v1961\(0) = '1' then
                \state\ <= q_wait1960;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$389\));
                \state\ <= pause_getI1958;
              end if;
            end if;
          when get_wait1971 =>
            if \$396_lock\(0) = '1' then
              \state\ <= get_wait1971;
            else
              \$395\ := \$396\;
              \$v1970\ := \$arr1451_ptr_take\;
              if \$v1970\(0) = '1' then
                \state\ <= q_wait1969;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$395\));
                \state\ <= pause_getI1967;
              end if;
            end if;
          when get_wait1976 =>
            if \$397_lock\(0) = '1' then
              \state\ <= get_wait1976;
            else
              \$381\ := \$397\;
              \$v1975\ := \$arr1452_ptr_take\;
              if \$v1975\(0) = '1' then
                \state\ <= q_wait1974;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1972;
              end if;
            end if;
          when get_wait1989 =>
            if \$418_lock\(0) = '1' then
              \state\ <= get_wait1989;
            else
              \$417\ := \$418\;
              \$v1988\ := \$arr1451_ptr_take\;
              if \$v1988\(0) = '1' then
                \state\ <= q_wait1987;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$417\));
                \state\ <= pause_getI1985;
              end if;
            end if;
          when get_wait1998 =>
            if \$424_lock\(0) = '1' then
              \state\ <= get_wait1998;
            else
              \$423\ := \$424\;
              \$v1997\ := \$arr1451_ptr_take\;
              if \$v1997\(0) = '1' then
                \state\ <= q_wait1996;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$423\));
                \state\ <= pause_getI1994;
              end if;
            end if;
          when get_wait2007 =>
            if \$433_lock\(0) = '1' then
              \state\ <= get_wait2007;
            else
              \$433_lock\ := eclat_true;
              \state\ <= get_pause2008;
            end if;
          when get_wait2009 =>
            if \$437_lock\(0) = '1' then
              \state\ <= get_wait2009;
            else
              \$436\ := \$437\;
              \$435\ := \$436\ & "00000000000000000000000000000001";
              \$434\ := eclat_sub(\$435\);
              if \$433_lock\(0) = '1' then
                \state\ <= get_wait2007;
              else
                \$433_lock\ := eclat_true;
                \state\ <= get_pause2008;
              end if;
            end if;
          when get_wait2024 =>
            if \$432_lock\(0) = '1' then
              \state\ <= get_wait2024;
            else
              \$432_lock\ := eclat_true;
              \state\ <= get_pause2025;
            end if;
          when get_wait2037 =>
            if \$438_lock\(0) = '1' then
              \state\ <= get_wait2037;
            else
              \$428_i\ := \$438\;
              \$v2036\ := eclat_gt(\$428_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2036\(0) = '1' then
                \$v2035\ := eclat_eq(\$428_i\ & X"000" & X"15f90");
                if \$v2035\(0) = '1' then
                  \$v2023\ := \$arr1451_ptr_take\;
                  if \$v2023\(0) = '1' then
                    \state\ <= q_wait2022;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2018\ := "00000000000000000000000000000000";
                    \$v2019\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$427_result_after_f\ & "0001" & \$v2018\ & "0001" & \$v2019\;
                    \state\ <= pause_setI2020;
                  end if;
                else
                  \$v2034\ := \$arr1451_ptr_take\;
                  if \$v2034\(0) = '1' then
                    \state\ <= q_wait2033;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2030\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$427_result_after_f\ & "0010" & \$428_i\ & "0001" & \$v2030\;
                    \state\ <= pause_setI2031;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811403\;
              end if;
            end if;
          when get_wait2049 =>
            if \$461_lock\(0) = '1' then
              \state\ <= get_wait2049;
            else
              \$461_lock\ := eclat_true;
              \state\ <= get_pause2050;
            end if;
          when get_wait2058 =>
            if \$473_lock\(0) = '1' then
              \state\ <= get_wait2058;
            else
              \$472\ := \$473\;
              \$v2057\ := \$arr1451_ptr_take\;
              if \$v2057\(0) = '1' then
                \state\ <= q_wait2056;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$472\));
                \state\ <= pause_getI2054;
              end if;
            end if;
          when get_wait2076 =>
            if \$453_lock\(0) = '1' then
              \state\ <= get_wait2076;
            else
              \$452\ := \$453\;
              \$v2075\ := \$arr1451_ptr_take\;
              if \$v2075\(0) = '1' then
                \state\ <= q_wait2074;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$452\));
                \state\ <= pause_getI2072;
              end if;
            end if;
          when get_wait2085 =>
            if \$459_lock\(0) = '1' then
              \state\ <= get_wait2085;
            else
              \$458\ := \$459\;
              \$v2084\ := \$arr1451_ptr_take\;
              if \$v2084\(0) = '1' then
                \state\ <= q_wait2083;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$458\));
                \state\ <= pause_getI2081;
              end if;
            end if;
          when get_wait2090 =>
            if \$460_lock\(0) = '1' then
              \state\ <= get_wait2090;
            else
              \$444\ := \$460\;
              \$v2089\ := \$arr1452_ptr_take\;
              if \$v2089\(0) = '1' then
                \state\ <= q_wait2088;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2086;
              end if;
            end if;
          when get_wait2103 =>
            if \$481_lock\(0) = '1' then
              \state\ <= get_wait2103;
            else
              \$480\ := \$481\;
              \$v2102\ := \$arr1451_ptr_take\;
              if \$v2102\(0) = '1' then
                \state\ <= q_wait2101;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$480\));
                \state\ <= pause_getI2099;
              end if;
            end if;
          when get_wait2112 =>
            if \$487_lock\(0) = '1' then
              \state\ <= get_wait2112;
            else
              \$486\ := \$487\;
              \$v2111\ := \$arr1451_ptr_take\;
              if \$v2111\(0) = '1' then
                \state\ <= q_wait2110;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$486\));
                \state\ <= pause_getI2108;
              end if;
            end if;
          when get_wait2117 =>
            if \$507_lock\(0) = '1' then
              \state\ <= get_wait2117;
            else
              \$507_lock\ := eclat_true;
              \state\ <= get_pause2118;
            end if;
          when get_wait2126 =>
            if \$519_lock\(0) = '1' then
              \state\ <= get_wait2126;
            else
              \$518\ := \$519\;
              \$v2125\ := \$arr1451_ptr_take\;
              if \$v2125\(0) = '1' then
                \state\ <= q_wait2124;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$518\));
                \state\ <= pause_getI2122;
              end if;
            end if;
          when get_wait2144 =>
            if \$499_lock\(0) = '1' then
              \state\ <= get_wait2144;
            else
              \$498\ := \$499\;
              \$v2143\ := \$arr1451_ptr_take\;
              if \$v2143\(0) = '1' then
                \state\ <= q_wait2142;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$498\));
                \state\ <= pause_getI2140;
              end if;
            end if;
          when get_wait2153 =>
            if \$505_lock\(0) = '1' then
              \state\ <= get_wait2153;
            else
              \$504\ := \$505\;
              \$v2152\ := \$arr1451_ptr_take\;
              if \$v2152\(0) = '1' then
                \state\ <= q_wait2151;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$504\));
                \state\ <= pause_getI2149;
              end if;
            end if;
          when get_wait2158 =>
            if \$506_lock\(0) = '1' then
              \state\ <= get_wait2158;
            else
              \$490\ := \$506\;
              \$v2157\ := \$arr1452_ptr_take\;
              if \$v2157\(0) = '1' then
                \state\ <= q_wait2156;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2154;
              end if;
            end if;
          when get_wait2171 =>
            if \$527_lock\(0) = '1' then
              \state\ <= get_wait2171;
            else
              \$526\ := \$527\;
              \$v2170\ := \$arr1451_ptr_take\;
              if \$v2170\(0) = '1' then
                \state\ <= q_wait2169;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$526\));
                \state\ <= pause_getI2167;
              end if;
            end if;
          when get_wait2180 =>
            if \$533_lock\(0) = '1' then
              \state\ <= get_wait2180;
            else
              \$532\ := \$533\;
              \$v2179\ := \$arr1451_ptr_take\;
              if \$v2179\(0) = '1' then
                \state\ <= q_wait2178;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$532\));
                \state\ <= pause_getI2176;
              end if;
            end if;
          when get_wait2189 =>
            if \$v58_lock\(0) = '1' then
              \state\ <= get_wait2189;
            else
              \$v58_lock\ := eclat_true;
              \state\ <= get_pause2190;
            end if;
          when get_wait2205 =>
            if \$v55_lock\(0) = '1' then
              \state\ <= get_wait2205;
            else
              \$v55_lock\ := eclat_true;
              \state\ <= get_pause2206;
            end if;
          when get_wait2229 =>
            if \$v45_lock\(0) = '1' then
              \state\ <= get_wait2229;
            else
              \$82_i\ := \$v45\;
              \$v2228\ := eclat_gt(\$82_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2228\(0) = '1' then
                \$v2227\ := eclat_eq(\$82_i\ & X"000" & X"15f90");
                if \$v2227\(0) = '1' then
                  \$v2204\ := \$arr1451_ptr_take\;
                  if \$v2204\(0) = '1' then
                    \state\ <= q_wait2203;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2198\ := "00000000000000000000000000000000";
                    \$v2199\ := "00000000000000000000000000000000";
                    \$v2200\ := "00000000000000000000000000000101";
                    \$v2195\ := "00000000000000000000000000000000";
                    \$v2196\ := "00000000000000000000000000000000";
                    \$v2197\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(result & "0001" & \$v2198\ & "0001" & \$v2199\ & "0001" & \$v2200\ & "0001" & \$v2195\ & "0001" & \$v2196\ & "0001" & \$v2197\);
                    \state\ <= pause_setI2201;
                  end if;
                else
                  \$v2226\ := \$arr1451_ptr_take\;
                  if \$v2226\(0) = '1' then
                    \state\ <= q_wait2225;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2220\ := "00000000000000000000000000000000";
                    \$v2221\ := "00000000000000000000000000000000";
                    \$v2222\ := "00000000000000000000000000000101";
                    \$v2217\ := "00000000000000000000000000000000";
                    \$v2218\ := "00000000000000000000000000000000";
                    \$v2219\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(result & "0001" & \$v2220\ & "0001" & \$v2221\ & "0001" & \$v2222\ & "0001" & \$v2217\ & "0001" & \$v2218\ & "0001" & \$v2219\);
                    \state\ <= pause_setI2223;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811408\;
              end if;
            end if;
          when get_wait2240 =>
            if \$559_lock\(0) = '1' then
              \state\ <= get_wait2240;
            else
              \$559_lock\ := eclat_true;
              \state\ <= get_pause2241;
            end if;
          when get_wait2249 =>
            if \$571_lock\(0) = '1' then
              \state\ <= get_wait2249;
            else
              \$570\ := \$571\;
              \$v2248\ := \$arr1451_ptr_take\;
              if \$v2248\(0) = '1' then
                \state\ <= q_wait2247;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$570\));
                \state\ <= pause_getI2245;
              end if;
            end if;
          when get_wait2267 =>
            if \$551_lock\(0) = '1' then
              \state\ <= get_wait2267;
            else
              \$550\ := \$551\;
              \$v2266\ := \$arr1451_ptr_take\;
              if \$v2266\(0) = '1' then
                \state\ <= q_wait2265;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$550\));
                \state\ <= pause_getI2263;
              end if;
            end if;
          when get_wait2276 =>
            if \$557_lock\(0) = '1' then
              \state\ <= get_wait2276;
            else
              \$556\ := \$557\;
              \$v2275\ := \$arr1451_ptr_take\;
              if \$v2275\(0) = '1' then
                \state\ <= q_wait2274;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$556\));
                \state\ <= pause_getI2272;
              end if;
            end if;
          when get_wait2281 =>
            if \$558_lock\(0) = '1' then
              \state\ <= get_wait2281;
            else
              \$542\ := \$558\;
              \$v2280\ := \$arr1452_ptr_take\;
              if \$v2280\(0) = '1' then
                \state\ <= q_wait2279;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2277;
              end if;
            end if;
          when get_wait2294 =>
            if \$579_lock\(0) = '1' then
              \state\ <= get_wait2294;
            else
              \$578\ := \$579\;
              \$v2293\ := \$arr1451_ptr_take\;
              if \$v2293\(0) = '1' then
                \state\ <= q_wait2292;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$578\));
                \state\ <= pause_getI2290;
              end if;
            end if;
          when get_wait2303 =>
            if \$585_lock\(0) = '1' then
              \state\ <= get_wait2303;
            else
              \$584\ := \$585\;
              \$v2302\ := \$arr1451_ptr_take\;
              if \$v2302\(0) = '1' then
                \state\ <= q_wait2301;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$584\));
                \state\ <= pause_getI2299;
              end if;
            end if;
          when get_wait2308 =>
            if \$605_lock\(0) = '1' then
              \state\ <= get_wait2308;
            else
              \$605_lock\ := eclat_true;
              \state\ <= get_pause2309;
            end if;
          when get_wait2317 =>
            if \$617_lock\(0) = '1' then
              \state\ <= get_wait2317;
            else
              \$616\ := \$617\;
              \$v2316\ := \$arr1451_ptr_take\;
              if \$v2316\(0) = '1' then
                \state\ <= q_wait2315;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$616\));
                \state\ <= pause_getI2313;
              end if;
            end if;
          when get_wait2335 =>
            if \$597_lock\(0) = '1' then
              \state\ <= get_wait2335;
            else
              \$596\ := \$597\;
              \$v2334\ := \$arr1451_ptr_take\;
              if \$v2334\(0) = '1' then
                \state\ <= q_wait2333;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$596\));
                \state\ <= pause_getI2331;
              end if;
            end if;
          when get_wait2344 =>
            if \$603_lock\(0) = '1' then
              \state\ <= get_wait2344;
            else
              \$602\ := \$603\;
              \$v2343\ := \$arr1451_ptr_take\;
              if \$v2343\(0) = '1' then
                \state\ <= q_wait2342;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$602\));
                \state\ <= pause_getI2340;
              end if;
            end if;
          when get_wait2349 =>
            if \$604_lock\(0) = '1' then
              \state\ <= get_wait2349;
            else
              \$588\ := \$604\;
              \$v2348\ := \$arr1452_ptr_take\;
              if \$v2348\(0) = '1' then
                \state\ <= q_wait2347;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2345;
              end if;
            end if;
          when get_wait2362 =>
            if \$625_lock\(0) = '1' then
              \state\ <= get_wait2362;
            else
              \$624\ := \$625\;
              \$v2361\ := \$arr1451_ptr_take\;
              if \$v2361\(0) = '1' then
                \state\ <= q_wait2360;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$624\));
                \state\ <= pause_getI2358;
              end if;
            end if;
          when get_wait2371 =>
            if \$631_lock\(0) = '1' then
              \state\ <= get_wait2371;
            else
              \$630\ := \$631\;
              \$v2370\ := \$arr1451_ptr_take\;
              if \$v2370\(0) = '1' then
                \state\ <= q_wait2369;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$630\));
                \state\ <= pause_getI2367;
              end if;
            end if;
          when get_wait2380 =>
            if \$640_lock\(0) = '1' then
              \state\ <= get_wait2380;
            else
              \$640_lock\ := eclat_true;
              \state\ <= get_pause2381;
            end if;
          when get_wait2396 =>
            if \$639_lock\(0) = '1' then
              \state\ <= get_wait2396;
            else
              \$639_lock\ := eclat_true;
              \state\ <= get_pause2397;
            end if;
          when get_wait2420 =>
            if \$641_lock\(0) = '1' then
              \state\ <= get_wait2420;
            else
              \$635_i\ := \$641\;
              \$v2419\ := eclat_gt(\$635_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2419\(0) = '1' then
                \$v2418\ := eclat_eq(\$635_i\ & X"000" & X"15f90");
                if \$v2418\(0) = '1' then
                  \$v2395\ := \$arr1451_ptr_take\;
                  if \$v2395\(0) = '1' then
                    \state\ <= q_wait2394;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2389\ := "00000000000000000000000000000000";
                    \$v2390\ := "00000000000000000000000000000000";
                    \$v2391\ := "00000000000000000000000000000101";
                    \$v2386\ := "00000000000000000000000000000000";
                    \$v2387\ := "00000000000000000000000000000000";
                    \$v2388\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2389\ & "0001" & \$v2390\ & "0001" & \$v2391\ & "0001" & \$v2386\ & "0001" & \$v2387\ & "0001" & \$v2388\);
                    \state\ <= pause_setI2392;
                  end if;
                else
                  \$v2417\ := \$arr1451_ptr_take\;
                  if \$v2417\(0) = '1' then
                    \state\ <= q_wait2416;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2411\ := "00000000000000000000000000000000";
                    \$v2412\ := "00000000000000000000000000000000";
                    \$v2413\ := "00000000000000000000000000000101";
                    \$v2408\ := "00000000000000000000000000000000";
                    \$v2409\ := "00000000000000000000000000000000";
                    \$v2410\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2411\ & "0001" & \$v2412\ & "0001" & \$v2413\ & "0001" & \$v2408\ & "0001" & \$v2409\ & "0001" & \$v2410\);
                    \state\ <= pause_setI2414;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811413\;
              end if;
            end if;
          when get_wait2434 =>
            if \$661_lock\(0) = '1' then
              \state\ <= get_wait2434;
            else
              \$661_lock\ := eclat_true;
              \state\ <= get_pause2435;
            end if;
          when get_wait2443 =>
            if \$673_lock\(0) = '1' then
              \state\ <= get_wait2443;
            else
              \$672\ := \$673\;
              \$v2442\ := \$arr1451_ptr_take\;
              if \$v2442\(0) = '1' then
                \state\ <= q_wait2441;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$672\));
                \state\ <= pause_getI2439;
              end if;
            end if;
          when get_wait2461 =>
            if \$653_lock\(0) = '1' then
              \state\ <= get_wait2461;
            else
              \$652\ := \$653\;
              \$v2460\ := \$arr1451_ptr_take\;
              if \$v2460\(0) = '1' then
                \state\ <= q_wait2459;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$652\));
                \state\ <= pause_getI2457;
              end if;
            end if;
          when get_wait2470 =>
            if \$659_lock\(0) = '1' then
              \state\ <= get_wait2470;
            else
              \$658\ := \$659\;
              \$v2469\ := \$arr1451_ptr_take\;
              if \$v2469\(0) = '1' then
                \state\ <= q_wait2468;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$658\));
                \state\ <= pause_getI2466;
              end if;
            end if;
          when get_wait2475 =>
            if \$660_lock\(0) = '1' then
              \state\ <= get_wait2475;
            else
              \$644\ := \$660\;
              \$v2474\ := \$arr1452_ptr_take\;
              if \$v2474\(0) = '1' then
                \state\ <= q_wait2473;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2471;
              end if;
            end if;
          when get_wait2488 =>
            if \$681_lock\(0) = '1' then
              \state\ <= get_wait2488;
            else
              \$680\ := \$681\;
              \$v2487\ := \$arr1451_ptr_take\;
              if \$v2487\(0) = '1' then
                \state\ <= q_wait2486;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$680\));
                \state\ <= pause_getI2484;
              end if;
            end if;
          when get_wait2497 =>
            if \$687_lock\(0) = '1' then
              \state\ <= get_wait2497;
            else
              \$686\ := \$687\;
              \$v2496\ := \$arr1451_ptr_take\;
              if \$v2496\(0) = '1' then
                \state\ <= q_wait2495;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$686\));
                \state\ <= pause_getI2493;
              end if;
            end if;
          when get_wait2502 =>
            if \$707_lock\(0) = '1' then
              \state\ <= get_wait2502;
            else
              \$707_lock\ := eclat_true;
              \state\ <= get_pause2503;
            end if;
          when get_wait2511 =>
            if \$719_lock\(0) = '1' then
              \state\ <= get_wait2511;
            else
              \$718\ := \$719\;
              \$v2510\ := \$arr1451_ptr_take\;
              if \$v2510\(0) = '1' then
                \state\ <= q_wait2509;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$718\));
                \state\ <= pause_getI2507;
              end if;
            end if;
          when get_wait2529 =>
            if \$699_lock\(0) = '1' then
              \state\ <= get_wait2529;
            else
              \$698\ := \$699\;
              \$v2528\ := \$arr1451_ptr_take\;
              if \$v2528\(0) = '1' then
                \state\ <= q_wait2527;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$698\));
                \state\ <= pause_getI2525;
              end if;
            end if;
          when get_wait2538 =>
            if \$705_lock\(0) = '1' then
              \state\ <= get_wait2538;
            else
              \$704\ := \$705\;
              \$v2537\ := \$arr1451_ptr_take\;
              if \$v2537\(0) = '1' then
                \state\ <= q_wait2536;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$704\));
                \state\ <= pause_getI2534;
              end if;
            end if;
          when get_wait2543 =>
            if \$706_lock\(0) = '1' then
              \state\ <= get_wait2543;
            else
              \$690\ := \$706\;
              \$v2542\ := \$arr1452_ptr_take\;
              if \$v2542\(0) = '1' then
                \state\ <= q_wait2541;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2539;
              end if;
            end if;
          when get_wait2556 =>
            if \$727_lock\(0) = '1' then
              \state\ <= get_wait2556;
            else
              \$726\ := \$727\;
              \$v2555\ := \$arr1451_ptr_take\;
              if \$v2555\(0) = '1' then
                \state\ <= q_wait2554;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$726\));
                \state\ <= pause_getI2552;
              end if;
            end if;
          when get_wait2565 =>
            if \$733_lock\(0) = '1' then
              \state\ <= get_wait2565;
            else
              \$732\ := \$733\;
              \$v2564\ := \$arr1451_ptr_take\;
              if \$v2564\(0) = '1' then
                \state\ <= q_wait2563;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$732\));
                \state\ <= pause_getI2561;
              end if;
            end if;
          when get_wait2574 =>
            if \$739_lock\(0) = '1' then
              \state\ <= get_wait2574;
            else
              \$739_lock\ := eclat_true;
              \state\ <= get_pause2575;
            end if;
          when get_wait2584 =>
            if \$738_lock\(0) = '1' then
              \state\ <= get_wait2584;
            else
              \$738_lock\ := eclat_true;
              \state\ <= get_pause2585;
            end if;
          when get_wait2602 =>
            if \$743_lock\(0) = '1' then
              \state\ <= get_wait2602;
            else
              \$734_i\ := \$743\;
              \$v2601\ := eclat_gt(\$734_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2601\(0) = '1' then
                \$v2600\ := eclat_eq(\$734_i\ & X"000" & X"15f90");
                if \$v2600\(0) = '1' then
                  \$v2583\ := \$arr1451_ptr_take\;
                  if \$v2583\(0) = '1' then
                    \state\ <= q_wait2582;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
                    \state\ <= pause_setI2580;
                  end if;
                else
                  \$v2599\ := \$arr1451_ptr_take\;
                  if \$v2599\(0) = '1' then
                    \state\ <= q_wait2598;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
                    \state\ <= pause_setI2596;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811416\;
              end if;
            end if;
          when get_wait2614 =>
            if \$766_lock\(0) = '1' then
              \state\ <= get_wait2614;
            else
              \$766_lock\ := eclat_true;
              \state\ <= get_pause2615;
            end if;
          when get_wait2623 =>
            if \$778_lock\(0) = '1' then
              \state\ <= get_wait2623;
            else
              \$777\ := \$778\;
              \$v2622\ := \$arr1451_ptr_take\;
              if \$v2622\(0) = '1' then
                \state\ <= q_wait2621;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$777\));
                \state\ <= pause_getI2619;
              end if;
            end if;
          when get_wait2641 =>
            if \$758_lock\(0) = '1' then
              \state\ <= get_wait2641;
            else
              \$757\ := \$758\;
              \$v2640\ := \$arr1451_ptr_take\;
              if \$v2640\(0) = '1' then
                \state\ <= q_wait2639;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$757\));
                \state\ <= pause_getI2637;
              end if;
            end if;
          when get_wait2650 =>
            if \$764_lock\(0) = '1' then
              \state\ <= get_wait2650;
            else
              \$763\ := \$764\;
              \$v2649\ := \$arr1451_ptr_take\;
              if \$v2649\(0) = '1' then
                \state\ <= q_wait2648;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$763\));
                \state\ <= pause_getI2646;
              end if;
            end if;
          when get_wait2655 =>
            if \$765_lock\(0) = '1' then
              \state\ <= get_wait2655;
            else
              \$749\ := \$765\;
              \$v2654\ := \$arr1452_ptr_take\;
              if \$v2654\(0) = '1' then
                \state\ <= q_wait2653;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2651;
              end if;
            end if;
          when get_wait2668 =>
            if \$786_lock\(0) = '1' then
              \state\ <= get_wait2668;
            else
              \$785\ := \$786\;
              \$v2667\ := \$arr1451_ptr_take\;
              if \$v2667\(0) = '1' then
                \state\ <= q_wait2666;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$785\));
                \state\ <= pause_getI2664;
              end if;
            end if;
          when get_wait2677 =>
            if \$792_lock\(0) = '1' then
              \state\ <= get_wait2677;
            else
              \$791\ := \$792\;
              \$v2676\ := \$arr1451_ptr_take\;
              if \$v2676\(0) = '1' then
                \state\ <= q_wait2675;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$791\));
                \state\ <= pause_getI2673;
              end if;
            end if;
          when get_wait2682 =>
            if \$812_lock\(0) = '1' then
              \state\ <= get_wait2682;
            else
              \$812_lock\ := eclat_true;
              \state\ <= get_pause2683;
            end if;
          when get_wait2691 =>
            if \$824_lock\(0) = '1' then
              \state\ <= get_wait2691;
            else
              \$823\ := \$824\;
              \$v2690\ := \$arr1451_ptr_take\;
              if \$v2690\(0) = '1' then
                \state\ <= q_wait2689;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$823\));
                \state\ <= pause_getI2687;
              end if;
            end if;
          when get_wait2709 =>
            if \$804_lock\(0) = '1' then
              \state\ <= get_wait2709;
            else
              \$803\ := \$804\;
              \$v2708\ := \$arr1451_ptr_take\;
              if \$v2708\(0) = '1' then
                \state\ <= q_wait2707;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$803\));
                \state\ <= pause_getI2705;
              end if;
            end if;
          when get_wait2718 =>
            if \$810_lock\(0) = '1' then
              \state\ <= get_wait2718;
            else
              \$809\ := \$810\;
              \$v2717\ := \$arr1451_ptr_take\;
              if \$v2717\(0) = '1' then
                \state\ <= q_wait2716;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$809\));
                \state\ <= pause_getI2714;
              end if;
            end if;
          when get_wait2723 =>
            if \$811_lock\(0) = '1' then
              \state\ <= get_wait2723;
            else
              \$795\ := \$811\;
              \$v2722\ := \$arr1452_ptr_take\;
              if \$v2722\(0) = '1' then
                \state\ <= q_wait2721;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2719;
              end if;
            end if;
          when get_wait2736 =>
            if \$832_lock\(0) = '1' then
              \state\ <= get_wait2736;
            else
              \$831\ := \$832\;
              \$v2735\ := \$arr1451_ptr_take\;
              if \$v2735\(0) = '1' then
                \state\ <= q_wait2734;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$831\));
                \state\ <= pause_getI2732;
              end if;
            end if;
          when get_wait2745 =>
            if \$838_lock\(0) = '1' then
              \state\ <= get_wait2745;
            else
              \$837\ := \$838\;
              \$v2744\ := \$arr1451_ptr_take\;
              if \$v2744\(0) = '1' then
                \state\ <= q_wait2743;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$837\));
                \state\ <= pause_getI2741;
              end if;
            end if;
          when get_wait2754 =>
            if \$846_lock\(0) = '1' then
              \state\ <= get_wait2754;
            else
              \$846_lock\ := eclat_true;
              \state\ <= get_pause2755;
            end if;
          when get_wait2764 =>
            if \$845_lock\(0) = '1' then
              \state\ <= get_wait2764;
            else
              \$845_lock\ := eclat_true;
              \state\ <= get_pause2765;
            end if;
          when get_wait2782 =>
            if \$850_lock\(0) = '1' then
              \state\ <= get_wait2782;
            else
              \$841_i\ := \$850\;
              \$v2781\ := eclat_gt(\$841_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2781\(0) = '1' then
                \$v2780\ := eclat_eq(\$841_i\ & X"000" & X"15f90");
                if \$v2780\(0) = '1' then
                  \$v2763\ := \$arr1451_ptr_take\;
                  if \$v2763\(0) = '1' then
                    \state\ <= q_wait2762;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
                    \state\ <= pause_setI2760;
                  end if;
                else
                  \$v2779\ := \$arr1451_ptr_take\;
                  if \$v2779\(0) = '1' then
                    \state\ <= q_wait2778;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
                    \state\ <= pause_setI2776;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811420\;
              end if;
            end if;
          when get_wait2794 =>
            if \$875_lock\(0) = '1' then
              \state\ <= get_wait2794;
            else
              \$875_lock\ := eclat_true;
              \state\ <= get_pause2795;
            end if;
          when get_wait2803 =>
            if \$887_lock\(0) = '1' then
              \state\ <= get_wait2803;
            else
              \$886\ := \$887\;
              \$v2802\ := \$arr1451_ptr_take\;
              if \$v2802\(0) = '1' then
                \state\ <= q_wait2801;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$886\));
                \state\ <= pause_getI2799;
              end if;
            end if;
          when get_wait2821 =>
            if \$867_lock\(0) = '1' then
              \state\ <= get_wait2821;
            else
              \$866\ := \$867\;
              \$v2820\ := \$arr1451_ptr_take\;
              if \$v2820\(0) = '1' then
                \state\ <= q_wait2819;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$866\));
                \state\ <= pause_getI2817;
              end if;
            end if;
          when get_wait2830 =>
            if \$873_lock\(0) = '1' then
              \state\ <= get_wait2830;
            else
              \$872\ := \$873\;
              \$v2829\ := \$arr1451_ptr_take\;
              if \$v2829\(0) = '1' then
                \state\ <= q_wait2828;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$872\));
                \state\ <= pause_getI2826;
              end if;
            end if;
          when get_wait2835 =>
            if \$874_lock\(0) = '1' then
              \state\ <= get_wait2835;
            else
              \$858\ := \$874\;
              \$v2834\ := \$arr1452_ptr_take\;
              if \$v2834\(0) = '1' then
                \state\ <= q_wait2833;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2831;
              end if;
            end if;
          when get_wait2848 =>
            if \$895_lock\(0) = '1' then
              \state\ <= get_wait2848;
            else
              \$894\ := \$895\;
              \$v2847\ := \$arr1451_ptr_take\;
              if \$v2847\(0) = '1' then
                \state\ <= q_wait2846;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$894\));
                \state\ <= pause_getI2844;
              end if;
            end if;
          when get_wait2857 =>
            if \$901_lock\(0) = '1' then
              \state\ <= get_wait2857;
            else
              \$900\ := \$901\;
              \$v2856\ := \$arr1451_ptr_take\;
              if \$v2856\(0) = '1' then
                \state\ <= q_wait2855;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$900\));
                \state\ <= pause_getI2853;
              end if;
            end if;
          when get_wait2862 =>
            if \$921_lock\(0) = '1' then
              \state\ <= get_wait2862;
            else
              \$921_lock\ := eclat_true;
              \state\ <= get_pause2863;
            end if;
          when get_wait2871 =>
            if \$933_lock\(0) = '1' then
              \state\ <= get_wait2871;
            else
              \$932\ := \$933\;
              \$v2870\ := \$arr1451_ptr_take\;
              if \$v2870\(0) = '1' then
                \state\ <= q_wait2869;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$932\));
                \state\ <= pause_getI2867;
              end if;
            end if;
          when get_wait2889 =>
            if \$913_lock\(0) = '1' then
              \state\ <= get_wait2889;
            else
              \$912\ := \$913\;
              \$v2888\ := \$arr1451_ptr_take\;
              if \$v2888\(0) = '1' then
                \state\ <= q_wait2887;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$912\));
                \state\ <= pause_getI2885;
              end if;
            end if;
          when get_wait2898 =>
            if \$919_lock\(0) = '1' then
              \state\ <= get_wait2898;
            else
              \$918\ := \$919\;
              \$v2897\ := \$arr1451_ptr_take\;
              if \$v2897\(0) = '1' then
                \state\ <= q_wait2896;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$918\));
                \state\ <= pause_getI2894;
              end if;
            end if;
          when get_wait2903 =>
            if \$920_lock\(0) = '1' then
              \state\ <= get_wait2903;
            else
              \$904\ := \$920\;
              \$v2902\ := \$arr1452_ptr_take\;
              if \$v2902\(0) = '1' then
                \state\ <= q_wait2901;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2899;
              end if;
            end if;
          when get_wait2916 =>
            if \$941_lock\(0) = '1' then
              \state\ <= get_wait2916;
            else
              \$940\ := \$941\;
              \$v2915\ := \$arr1451_ptr_take\;
              if \$v2915\(0) = '1' then
                \state\ <= q_wait2914;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$940\));
                \state\ <= pause_getI2912;
              end if;
            end if;
          when get_wait2925 =>
            if \$947_lock\(0) = '1' then
              \state\ <= get_wait2925;
            else
              \$946\ := \$947\;
              \$v2924\ := \$arr1451_ptr_take\;
              if \$v2924\(0) = '1' then
                \state\ <= q_wait2923;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$946\));
                \state\ <= pause_getI2921;
              end if;
            end if;
          when get_wait2934 =>
            if \$955_lock\(0) = '1' then
              \state\ <= get_wait2934;
            else
              \$955_lock\ := eclat_true;
              \state\ <= get_pause2935;
            end if;
          when get_wait2944 =>
            if \$954_lock\(0) = '1' then
              \state\ <= get_wait2944;
            else
              \$954_lock\ := eclat_true;
              \state\ <= get_pause2945;
            end if;
          when get_wait2962 =>
            if \$959_lock\(0) = '1' then
              \state\ <= get_wait2962;
            else
              \$950_i\ := \$959\;
              \$v2961\ := eclat_gt(\$950_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2961\(0) = '1' then
                \$v2960\ := eclat_eq(\$950_i\ & X"000" & X"15f90");
                if \$v2960\(0) = '1' then
                  \$v2943\ := \$arr1451_ptr_take\;
                  if \$v2943\(0) = '1' then
                    \state\ <= q_wait2942;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
                    \state\ <= pause_setI2940;
                  end if;
                else
                  \$v2959\ := \$arr1451_ptr_take\;
                  if \$v2959\(0) = '1' then
                    \state\ <= q_wait2958;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
                    \state\ <= pause_setI2956;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811424\;
              end if;
            end if;
          when get_wait2974 =>
            if \$984_lock\(0) = '1' then
              \state\ <= get_wait2974;
            else
              \$984_lock\ := eclat_true;
              \state\ <= get_pause2975;
            end if;
          when get_wait2983 =>
            if \$996_lock\(0) = '1' then
              \state\ <= get_wait2983;
            else
              \$995\ := \$996\;
              \$v2982\ := \$arr1451_ptr_take\;
              if \$v2982\(0) = '1' then
                \state\ <= q_wait2981;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$995\));
                \state\ <= pause_getI2979;
              end if;
            end if;
          when get_wait3001 =>
            if \$976_lock\(0) = '1' then
              \state\ <= get_wait3001;
            else
              \$975\ := \$976\;
              \$v3000\ := \$arr1451_ptr_take\;
              if \$v3000\(0) = '1' then
                \state\ <= q_wait2999;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$975\));
                \state\ <= pause_getI2997;
              end if;
            end if;
          when get_wait3010 =>
            if \$982_lock\(0) = '1' then
              \state\ <= get_wait3010;
            else
              \$981\ := \$982\;
              \$v3009\ := \$arr1451_ptr_take\;
              if \$v3009\(0) = '1' then
                \state\ <= q_wait3008;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$981\));
                \state\ <= pause_getI3006;
              end if;
            end if;
          when get_wait3015 =>
            if \$983_lock\(0) = '1' then
              \state\ <= get_wait3015;
            else
              \$967\ := \$983\;
              \$v3014\ := \$arr1452_ptr_take\;
              if \$v3014\(0) = '1' then
                \state\ <= q_wait3013;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3011;
              end if;
            end if;
          when get_wait3028 =>
            if \$1004_lock\(0) = '1' then
              \state\ <= get_wait3028;
            else
              \$1003\ := \$1004\;
              \$v3027\ := \$arr1451_ptr_take\;
              if \$v3027\(0) = '1' then
                \state\ <= q_wait3026;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1003\));
                \state\ <= pause_getI3024;
              end if;
            end if;
          when get_wait3037 =>
            if \$1010_lock\(0) = '1' then
              \state\ <= get_wait3037;
            else
              \$1009\ := \$1010\;
              \$v3036\ := \$arr1451_ptr_take\;
              if \$v3036\(0) = '1' then
                \state\ <= q_wait3035;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1009\));
                \state\ <= pause_getI3033;
              end if;
            end if;
          when get_wait3042 =>
            if \$1030_lock\(0) = '1' then
              \state\ <= get_wait3042;
            else
              \$1030_lock\ := eclat_true;
              \state\ <= get_pause3043;
            end if;
          when get_wait3051 =>
            if \$1042_lock\(0) = '1' then
              \state\ <= get_wait3051;
            else
              \$1041\ := \$1042\;
              \$v3050\ := \$arr1451_ptr_take\;
              if \$v3050\(0) = '1' then
                \state\ <= q_wait3049;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1041\));
                \state\ <= pause_getI3047;
              end if;
            end if;
          when get_wait3069 =>
            if \$1022_lock\(0) = '1' then
              \state\ <= get_wait3069;
            else
              \$1021\ := \$1022\;
              \$v3068\ := \$arr1451_ptr_take\;
              if \$v3068\(0) = '1' then
                \state\ <= q_wait3067;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1021\));
                \state\ <= pause_getI3065;
              end if;
            end if;
          when get_wait3078 =>
            if \$1028_lock\(0) = '1' then
              \state\ <= get_wait3078;
            else
              \$1027\ := \$1028\;
              \$v3077\ := \$arr1451_ptr_take\;
              if \$v3077\(0) = '1' then
                \state\ <= q_wait3076;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1027\));
                \state\ <= pause_getI3074;
              end if;
            end if;
          when get_wait3083 =>
            if \$1029_lock\(0) = '1' then
              \state\ <= get_wait3083;
            else
              \$1013\ := \$1029\;
              \$v3082\ := \$arr1452_ptr_take\;
              if \$v3082\(0) = '1' then
                \state\ <= q_wait3081;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3079;
              end if;
            end if;
          when get_wait3096 =>
            if \$1050_lock\(0) = '1' then
              \state\ <= get_wait3096;
            else
              \$1049\ := \$1050\;
              \$v3095\ := \$arr1451_ptr_take\;
              if \$v3095\(0) = '1' then
                \state\ <= q_wait3094;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1049\));
                \state\ <= pause_getI3092;
              end if;
            end if;
          when get_wait3105 =>
            if \$1056_lock\(0) = '1' then
              \state\ <= get_wait3105;
            else
              \$1055\ := \$1056\;
              \$v3104\ := \$arr1451_ptr_take\;
              if \$v3104\(0) = '1' then
                \state\ <= q_wait3103;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1055\));
                \state\ <= pause_getI3101;
              end if;
            end if;
          when get_wait3114 =>
            if \$1065_lock\(0) = '1' then
              \state\ <= get_wait3114;
            else
              \$1065_lock\ := eclat_true;
              \state\ <= get_pause3115;
            end if;
          when get_wait3116 =>
            if \$1069_lock\(0) = '1' then
              \state\ <= get_wait3116;
            else
              \$1068\ := \$1069\;
              \$1067\ := \$1068\ & "00000000000000000000000000000001";
              \$1066\ := eclat_sub(\$1067\);
              if \$1065_lock\(0) = '1' then
                \state\ <= get_wait3114;
              else
                \$1065_lock\ := eclat_true;
                \state\ <= get_pause3115;
              end if;
            end if;
          when get_wait3131 =>
            if \$1061_lock\(0) = '1' then
              \state\ <= get_wait3131;
            else
              \$1061_lock\ := eclat_true;
              \state\ <= get_pause3132;
            end if;
          when get_wait3144 =>
            if \$1073_lock\(0) = '1' then
              \state\ <= get_wait3144;
            else
              \$1057_i\ := \$1073\;
              \$v3143\ := eclat_gt(\$1057_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3143\(0) = '1' then
                \$v3142\ := eclat_eq(\$1057_i\ & X"000" & X"15f90");
                if \$v3142\(0) = '1' then
                  \$v3130\ := \$arr1451_ptr_take\;
                  if \$v3130\(0) = '1' then
                    \state\ <= q_wait3129;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3125\ := "00000000000000000000000000000000";
                    \$v3126\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$58_result\(72 to 107) & "0001" & \$v3125\ & "0001" & \$v3126\;
                    \state\ <= pause_setI3127;
                  end if;
                else
                  \$v3141\ := \$arr1451_ptr_take\;
                  if \$v3141\(0) = '1' then
                    \state\ <= q_wait3140;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3137\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$58_result\(72 to 107) & "0010" & \$1057_i\ & "0001" & \$v3137\;
                    \state\ <= pause_setI3138;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811428\;
              end if;
            end if;
          when get_wait3156 =>
            if \$1098_lock\(0) = '1' then
              \state\ <= get_wait3156;
            else
              \$1098_lock\ := eclat_true;
              \state\ <= get_pause3157;
            end if;
          when get_wait3165 =>
            if \$1110_lock\(0) = '1' then
              \state\ <= get_wait3165;
            else
              \$1109\ := \$1110\;
              \$v3164\ := \$arr1451_ptr_take\;
              if \$v3164\(0) = '1' then
                \state\ <= q_wait3163;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1109\));
                \state\ <= pause_getI3161;
              end if;
            end if;
          when get_wait3183 =>
            if \$1090_lock\(0) = '1' then
              \state\ <= get_wait3183;
            else
              \$1089\ := \$1090\;
              \$v3182\ := \$arr1451_ptr_take\;
              if \$v3182\(0) = '1' then
                \state\ <= q_wait3181;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1089\));
                \state\ <= pause_getI3179;
              end if;
            end if;
          when get_wait3192 =>
            if \$1096_lock\(0) = '1' then
              \state\ <= get_wait3192;
            else
              \$1095\ := \$1096\;
              \$v3191\ := \$arr1451_ptr_take\;
              if \$v3191\(0) = '1' then
                \state\ <= q_wait3190;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1095\));
                \state\ <= pause_getI3188;
              end if;
            end if;
          when get_wait3197 =>
            if \$1097_lock\(0) = '1' then
              \state\ <= get_wait3197;
            else
              \$1081\ := \$1097\;
              \$v3196\ := \$arr1452_ptr_take\;
              if \$v3196\(0) = '1' then
                \state\ <= q_wait3195;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3193;
              end if;
            end if;
          when get_wait3210 =>
            if \$1118_lock\(0) = '1' then
              \state\ <= get_wait3210;
            else
              \$1117\ := \$1118\;
              \$v3209\ := \$arr1451_ptr_take\;
              if \$v3209\(0) = '1' then
                \state\ <= q_wait3208;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1117\));
                \state\ <= pause_getI3206;
              end if;
            end if;
          when get_wait3219 =>
            if \$1124_lock\(0) = '1' then
              \state\ <= get_wait3219;
            else
              \$1123\ := \$1124\;
              \$v3218\ := \$arr1451_ptr_take\;
              if \$v3218\(0) = '1' then
                \state\ <= q_wait3217;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1123\));
                \state\ <= pause_getI3215;
              end if;
            end if;
          when get_wait3228 =>
            if \$1134_lock\(0) = '1' then
              \state\ <= get_wait3228;
            else
              \$1134_lock\ := eclat_true;
              \state\ <= get_pause3229;
            end if;
          when get_wait3230 =>
            if \$1138_lock\(0) = '1' then
              \state\ <= get_wait3230;
            else
              \$1137\ := \$1138\;
              \$1136\ := \$1137\ & "00000000000000000000000000000001";
              \$1135\ := eclat_sub(\$1136\);
              if \$1134_lock\(0) = '1' then
                \state\ <= get_wait3228;
              else
                \$1134_lock\ := eclat_true;
                \state\ <= get_pause3229;
              end if;
            end if;
          when get_wait3245 =>
            if \$1130_lock\(0) = '1' then
              \state\ <= get_wait3245;
            else
              \$1130_lock\ := eclat_true;
              \state\ <= get_pause3246;
            end if;
          when get_wait3258 =>
            if \$1142_lock\(0) = '1' then
              \state\ <= get_wait3258;
            else
              \$1126_i\ := \$1142\;
              \$v3257\ := eclat_gt(\$1126_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3257\(0) = '1' then
                \$v3256\ := eclat_eq(\$1126_i\ & X"000" & X"15f90");
                if \$v3256\(0) = '1' then
                  \$v3244\ := \$arr1451_ptr_take\;
                  if \$v3244\(0) = '1' then
                    \state\ <= q_wait3243;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3239\ := "00000000000000000000000000000000";
                    \$v3240\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1125_result\(36 to 71) & "0001" & \$v3239\ & "0001" & \$v3240\;
                    \state\ <= pause_setI3241;
                  end if;
                else
                  \$v3255\ := \$arr1451_ptr_take\;
                  if \$v3255\(0) = '1' then
                    \state\ <= q_wait3254;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3251\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1125_result\(36 to 71) & "0010" & \$1126_i\ & "0001" & \$v3251\;
                    \state\ <= pause_setI3252;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811431\;
              end if;
            end if;
          when get_wait3270 =>
            if \$1167_lock\(0) = '1' then
              \state\ <= get_wait3270;
            else
              \$1167_lock\ := eclat_true;
              \state\ <= get_pause3271;
            end if;
          when get_wait3279 =>
            if \$1179_lock\(0) = '1' then
              \state\ <= get_wait3279;
            else
              \$1178\ := \$1179\;
              \$v3278\ := \$arr1451_ptr_take\;
              if \$v3278\(0) = '1' then
                \state\ <= q_wait3277;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1178\));
                \state\ <= pause_getI3275;
              end if;
            end if;
          when get_wait3297 =>
            if \$1159_lock\(0) = '1' then
              \state\ <= get_wait3297;
            else
              \$1158\ := \$1159\;
              \$v3296\ := \$arr1451_ptr_take\;
              if \$v3296\(0) = '1' then
                \state\ <= q_wait3295;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1158\));
                \state\ <= pause_getI3293;
              end if;
            end if;
          when get_wait3306 =>
            if \$1165_lock\(0) = '1' then
              \state\ <= get_wait3306;
            else
              \$1164\ := \$1165\;
              \$v3305\ := \$arr1451_ptr_take\;
              if \$v3305\(0) = '1' then
                \state\ <= q_wait3304;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1164\));
                \state\ <= pause_getI3302;
              end if;
            end if;
          when get_wait3311 =>
            if \$1166_lock\(0) = '1' then
              \state\ <= get_wait3311;
            else
              \$1150\ := \$1166\;
              \$v3310\ := \$arr1452_ptr_take\;
              if \$v3310\(0) = '1' then
                \state\ <= q_wait3309;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3307;
              end if;
            end if;
          when get_wait3324 =>
            if \$1187_lock\(0) = '1' then
              \state\ <= get_wait3324;
            else
              \$1186\ := \$1187\;
              \$v3323\ := \$arr1451_ptr_take\;
              if \$v3323\(0) = '1' then
                \state\ <= q_wait3322;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1186\));
                \state\ <= pause_getI3320;
              end if;
            end if;
          when get_wait3333 =>
            if \$1193_lock\(0) = '1' then
              \state\ <= get_wait3333;
            else
              \$1192\ := \$1193\;
              \$v3332\ := \$arr1451_ptr_take\;
              if \$v3332\(0) = '1' then
                \state\ <= q_wait3331;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1192\));
                \state\ <= pause_getI3329;
              end if;
            end if;
          when get_wait3342 =>
            if \$1203_lock\(0) = '1' then
              \state\ <= get_wait3342;
            else
              \$1203_lock\ := eclat_true;
              \state\ <= get_pause3343;
            end if;
          when get_wait3344 =>
            if \$1207_lock\(0) = '1' then
              \state\ <= get_wait3344;
            else
              \$1206\ := \$1207\;
              \$1205\ := \$1206\ & "00000000000000000000000000000001";
              \$1204\ := eclat_sub(\$1205\);
              if \$1203_lock\(0) = '1' then
                \state\ <= get_wait3342;
              else
                \$1203_lock\ := eclat_true;
                \state\ <= get_pause3343;
              end if;
            end if;
          when get_wait3359 =>
            if \$1199_lock\(0) = '1' then
              \state\ <= get_wait3359;
            else
              \$1199_lock\ := eclat_true;
              \state\ <= get_pause3360;
            end if;
          when get_wait3372 =>
            if \$1211_lock\(0) = '1' then
              \state\ <= get_wait3372;
            else
              \$1195_i\ := \$1211\;
              \$v3371\ := eclat_gt(\$1195_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3371\(0) = '1' then
                \$v3370\ := eclat_eq(\$1195_i\ & X"000" & X"15f90");
                if \$v3370\(0) = '1' then
                  \$v3358\ := \$arr1451_ptr_take\;
                  if \$v3358\(0) = '1' then
                    \state\ <= q_wait3357;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3353\ := "00000000000000000000000000000000";
                    \$v3354\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1194_result\(0 to 35) & "0001" & \$v3353\ & "0001" & \$v3354\;
                    \state\ <= pause_setI3355;
                  end if;
                else
                  \$v3369\ := \$arr1451_ptr_take\;
                  if \$v3369\(0) = '1' then
                    \state\ <= q_wait3368;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3365\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1194_result\(0 to 35) & "0010" & \$1195_i\ & "0001" & \$v3365\;
                    \state\ <= pause_setI3366;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811434\;
              end if;
            end if;
          when get_wait3384 =>
            if \$1236_lock\(0) = '1' then
              \state\ <= get_wait3384;
            else
              \$1236_lock\ := eclat_true;
              \state\ <= get_pause3385;
            end if;
          when get_wait3393 =>
            if \$1248_lock\(0) = '1' then
              \state\ <= get_wait3393;
            else
              \$1247\ := \$1248\;
              \$v3392\ := \$arr1451_ptr_take\;
              if \$v3392\(0) = '1' then
                \state\ <= q_wait3391;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1247\));
                \state\ <= pause_getI3389;
              end if;
            end if;
          when get_wait3411 =>
            if \$1228_lock\(0) = '1' then
              \state\ <= get_wait3411;
            else
              \$1227\ := \$1228\;
              \$v3410\ := \$arr1451_ptr_take\;
              if \$v3410\(0) = '1' then
                \state\ <= q_wait3409;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1227\));
                \state\ <= pause_getI3407;
              end if;
            end if;
          when get_wait3420 =>
            if \$1234_lock\(0) = '1' then
              \state\ <= get_wait3420;
            else
              \$1233\ := \$1234\;
              \$v3419\ := \$arr1451_ptr_take\;
              if \$v3419\(0) = '1' then
                \state\ <= q_wait3418;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1233\));
                \state\ <= pause_getI3416;
              end if;
            end if;
          when get_wait3425 =>
            if \$1235_lock\(0) = '1' then
              \state\ <= get_wait3425;
            else
              \$1219\ := \$1235\;
              \$v3424\ := \$arr1452_ptr_take\;
              if \$v3424\(0) = '1' then
                \state\ <= q_wait3423;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3421;
              end if;
            end if;
          when get_wait3438 =>
            if \$1256_lock\(0) = '1' then
              \state\ <= get_wait3438;
            else
              \$1255\ := \$1256\;
              \$v3437\ := \$arr1451_ptr_take\;
              if \$v3437\(0) = '1' then
                \state\ <= q_wait3436;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1255\));
                \state\ <= pause_getI3434;
              end if;
            end if;
          when get_wait3447 =>
            if \$1262_lock\(0) = '1' then
              \state\ <= get_wait3447;
            else
              \$1261\ := \$1262\;
              \$v3446\ := \$arr1451_ptr_take\;
              if \$v3446\(0) = '1' then
                \state\ <= q_wait3445;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1261\));
                \state\ <= pause_getI3443;
              end if;
            end if;
          when get_wait3456 =>
            if \$1268_lock\(0) = '1' then
              \state\ <= get_wait3456;
            else
              \$1268_lock\ := eclat_true;
              \state\ <= get_pause3457;
            end if;
          when get_wait3466 =>
            if \$1267_lock\(0) = '1' then
              \state\ <= get_wait3466;
            else
              \$1267_lock\ := eclat_true;
              \state\ <= get_pause3467;
            end if;
          when get_wait3484 =>
            if \$1269_lock\(0) = '1' then
              \state\ <= get_wait3484;
            else
              \$1263_i\ := \$1269\;
              \$v3483\ := eclat_gt(\$1263_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3483\(0) = '1' then
                \$v3482\ := eclat_eq(\$1263_i\ & X"000" & X"15f90");
                if \$v3482\(0) = '1' then
                  \$v3465\ := \$arr1451_ptr_take\;
                  if \$v3465\(0) = '1' then
                    \state\ <= q_wait3464;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$74_result_after_f\;
                    \state\ <= pause_setI3462;
                  end if;
                else
                  \$v3481\ := \$arr1451_ptr_take\;
                  if \$v3481\(0) = '1' then
                    \state\ <= q_wait3480;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$74_result_after_f\;
                    \state\ <= pause_setI3478;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811437\;
              end if;
            end if;
          when get_wait3498 =>
            if \$1289_lock\(0) = '1' then
              \state\ <= get_wait3498;
            else
              \$1289_lock\ := eclat_true;
              \state\ <= get_pause3499;
            end if;
          when get_wait3507 =>
            if \$1301_lock\(0) = '1' then
              \state\ <= get_wait3507;
            else
              \$1300\ := \$1301\;
              \$v3506\ := \$arr1451_ptr_take\;
              if \$v3506\(0) = '1' then
                \state\ <= q_wait3505;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1300\));
                \state\ <= pause_getI3503;
              end if;
            end if;
          when get_wait3525 =>
            if \$1281_lock\(0) = '1' then
              \state\ <= get_wait3525;
            else
              \$1280\ := \$1281\;
              \$v3524\ := \$arr1451_ptr_take\;
              if \$v3524\(0) = '1' then
                \state\ <= q_wait3523;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1280\));
                \state\ <= pause_getI3521;
              end if;
            end if;
          when get_wait3534 =>
            if \$1287_lock\(0) = '1' then
              \state\ <= get_wait3534;
            else
              \$1286\ := \$1287\;
              \$v3533\ := \$arr1451_ptr_take\;
              if \$v3533\(0) = '1' then
                \state\ <= q_wait3532;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1286\));
                \state\ <= pause_getI3530;
              end if;
            end if;
          when get_wait3539 =>
            if \$1288_lock\(0) = '1' then
              \state\ <= get_wait3539;
            else
              \$1272\ := \$1288\;
              \$v3538\ := \$arr1452_ptr_take\;
              if \$v3538\(0) = '1' then
                \state\ <= q_wait3537;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3535;
              end if;
            end if;
          when get_wait3552 =>
            if \$1309_lock\(0) = '1' then
              \state\ <= get_wait3552;
            else
              \$1308\ := \$1309\;
              \$v3551\ := \$arr1451_ptr_take\;
              if \$v3551\(0) = '1' then
                \state\ <= q_wait3550;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1308\));
                \state\ <= pause_getI3548;
              end if;
            end if;
          when get_wait3561 =>
            if \$1315_lock\(0) = '1' then
              \state\ <= get_wait3561;
            else
              \$1314\ := \$1315\;
              \$v3560\ := \$arr1451_ptr_take\;
              if \$v3560\(0) = '1' then
                \state\ <= q_wait3559;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1314\));
                \state\ <= pause_getI3557;
              end if;
            end if;
          when get_wait3570 =>
            if \$1324_lock\(0) = '1' then
              \state\ <= get_wait3570;
            else
              \$1324_lock\ := eclat_true;
              \state\ <= get_pause3571;
            end if;
          when get_wait3581 =>
            if \$1320_lock\(0) = '1' then
              \state\ <= get_wait3581;
            else
              \$1320_lock\ := eclat_true;
              \state\ <= get_pause3582;
            end if;
          when get_wait3600 =>
            if \$1328_lock\(0) = '1' then
              \state\ <= get_wait3600;
            else
              \$1316_i\ := \$1328\;
              \$v3599\ := eclat_gt(\$1316_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3599\(0) = '1' then
                \$v3598\ := eclat_eq(\$1316_i\ & X"000" & X"15f90");
                if \$v3598\(0) = '1' then
                  \$v3580\ := \$arr1451_ptr_take\;
                  if \$v3580\(0) = '1' then
                    \state\ <= q_wait3579;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3576\ := "00000000000000000000000000000001";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3576\;
                    \state\ <= pause_setI3577;
                  end if;
                else
                  \$v3597\ := \$arr1451_ptr_take\;
                  if \$v3597\(0) = '1' then
                    \state\ <= q_wait3596;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3593\ := "00000000000000000000000000000001";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3593\;
                    \state\ <= pause_setI3594;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811439\;
              end if;
            end if;
          when get_wait3609 =>
            if \$v78_lock\(0) = '1' then
              \state\ <= get_wait3609;
            else
              \$v79\ := \$v78\;
              \$v3608\ := \$arr1451_ptr_take\;
              if \$v3608\(0) = '1' then
                \state\ <= q_wait3607;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v79\));
                \state\ <= pause_getI3605;
              end if;
            end if;
          when get_wait3621 =>
            if \$1356_lock\(0) = '1' then
              \state\ <= get_wait3621;
            else
              \$1356_lock\ := eclat_true;
              \state\ <= get_pause3622;
            end if;
          when get_wait3630 =>
            if \$1368_lock\(0) = '1' then
              \state\ <= get_wait3630;
            else
              \$1367\ := \$1368\;
              \$v3629\ := \$arr1451_ptr_take\;
              if \$v3629\(0) = '1' then
                \state\ <= q_wait3628;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1367\));
                \state\ <= pause_getI3626;
              end if;
            end if;
          when get_wait3648 =>
            if \$1348_lock\(0) = '1' then
              \state\ <= get_wait3648;
            else
              \$1347\ := \$1348\;
              \$v3647\ := \$arr1451_ptr_take\;
              if \$v3647\(0) = '1' then
                \state\ <= q_wait3646;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1347\));
                \state\ <= pause_getI3644;
              end if;
            end if;
          when get_wait3657 =>
            if \$1354_lock\(0) = '1' then
              \state\ <= get_wait3657;
            else
              \$1353\ := \$1354\;
              \$v3656\ := \$arr1451_ptr_take\;
              if \$v3656\(0) = '1' then
                \state\ <= q_wait3655;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1353\));
                \state\ <= pause_getI3653;
              end if;
            end if;
          when get_wait3662 =>
            if \$1355_lock\(0) = '1' then
              \state\ <= get_wait3662;
            else
              \$1339\ := \$1355\;
              \$v3661\ := \$arr1452_ptr_take\;
              if \$v3661\(0) = '1' then
                \state\ <= q_wait3660;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3658;
              end if;
            end if;
          when get_wait3675 =>
            if \$1376_lock\(0) = '1' then
              \state\ <= get_wait3675;
            else
              \$1375\ := \$1376\;
              \$v3674\ := \$arr1451_ptr_take\;
              if \$v3674\(0) = '1' then
                \state\ <= q_wait3673;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1375\));
                \state\ <= pause_getI3671;
              end if;
            end if;
          when get_wait3684 =>
            if \$1382_lock\(0) = '1' then
              \state\ <= get_wait3684;
            else
              \$1381\ := \$1382\;
              \$v3683\ := \$arr1451_ptr_take\;
              if \$v3683\(0) = '1' then
                \state\ <= q_wait3682;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1381\));
                \state\ <= pause_getI3680;
              end if;
            end if;
          when get_wait3693 =>
            if \$1390_lock\(0) = '1' then
              \state\ <= get_wait3693;
            else
              \$1390_lock\ := eclat_true;
              \state\ <= get_pause3694;
            end if;
          when get_wait3695 =>
            if \$1394_lock\(0) = '1' then
              \state\ <= get_wait3695;
            else
              \$1393\ := \$1394\;
              \$1392\ := \$1393\ & "00000000000000000000000000000001";
              \$1391\ := eclat_sub(\$1392\);
              if \$1390_lock\(0) = '1' then
                \state\ <= get_wait3693;
              else
                \$1390_lock\ := eclat_true;
                \state\ <= get_pause3694;
              end if;
            end if;
          when get_wait3710 =>
            if \$1389_lock\(0) = '1' then
              \state\ <= get_wait3710;
            else
              \$1389_lock\ := eclat_true;
              \state\ <= get_pause3711;
            end if;
          when get_wait3723 =>
            if \$1395_lock\(0) = '1' then
              \state\ <= get_wait3723;
            else
              \$1385_i\ := \$1395\;
              \$v3722\ := eclat_gt(\$1385_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3722\(0) = '1' then
                \$v3721\ := eclat_eq(\$1385_i\ & X"000" & X"15f90");
                if \$v3721\(0) = '1' then
                  \$v3709\ := \$arr1451_ptr_take\;
                  if \$v3709\(0) = '1' then
                    \state\ <= q_wait3708;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3704\ := "00000000000000000000000000000000";
                    \$v3705\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1383_x\ & "0001" & \$v3704\ & "0001" & \$v3705\;
                    \state\ <= pause_setI3706;
                  end if;
                else
                  \$v3720\ := \$arr1451_ptr_take\;
                  if \$v3720\(0) = '1' then
                    \state\ <= q_wait3719;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3716\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1383_x\ & "0010" & \$1385_i\ & "0001" & \$v3716\;
                    \state\ <= pause_setI3717;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811442\;
              end if;
            end if;
          when get_wait3728 =>
            if \$1415_lock\(0) = '1' then
              \state\ <= get_wait3728;
            else
              \$1415_lock\ := eclat_true;
              \state\ <= get_pause3729;
            end if;
          when get_wait3737 =>
            if \$1427_lock\(0) = '1' then
              \state\ <= get_wait3737;
            else
              \$1426\ := \$1427\;
              \$v3736\ := \$arr1451_ptr_take\;
              if \$v3736\(0) = '1' then
                \state\ <= q_wait3735;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1426\));
                \state\ <= pause_getI3733;
              end if;
            end if;
          when get_wait3755 =>
            if \$1407_lock\(0) = '1' then
              \state\ <= get_wait3755;
            else
              \$1406\ := \$1407\;
              \$v3754\ := \$arr1451_ptr_take\;
              if \$v3754\(0) = '1' then
                \state\ <= q_wait3753;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1406\));
                \state\ <= pause_getI3751;
              end if;
            end if;
          when get_wait3764 =>
            if \$1413_lock\(0) = '1' then
              \state\ <= get_wait3764;
            else
              \$1412\ := \$1413\;
              \$v3763\ := \$arr1451_ptr_take\;
              if \$v3763\(0) = '1' then
                \state\ <= q_wait3762;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1412\));
                \state\ <= pause_getI3760;
              end if;
            end if;
          when get_wait3769 =>
            if \$1414_lock\(0) = '1' then
              \state\ <= get_wait3769;
            else
              \$1398\ := \$1414\;
              \$v3768\ := \$arr1452_ptr_take\;
              if \$v3768\(0) = '1' then
                \state\ <= q_wait3767;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3765;
              end if;
            end if;
          when get_wait3782 =>
            if \$1435_lock\(0) = '1' then
              \state\ <= get_wait3782;
            else
              \$1434\ := \$1435\;
              \$v3781\ := \$arr1451_ptr_take\;
              if \$v3781\(0) = '1' then
                \state\ <= q_wait3780;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1434\));
                \state\ <= pause_getI3778;
              end if;
            end if;
          when get_wait3791 =>
            if \$1441_lock\(0) = '1' then
              \state\ <= get_wait3791;
            else
              \$1440\ := \$1441\;
              \$v3790\ := \$arr1451_ptr_take\;
              if \$v3790\(0) = '1' then
                \state\ <= q_wait3789;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1440\));
                \state\ <= pause_getI3787;
              end if;
            end if;
          when get_wait3796 =>
            if \$1461_lock\(0) = '1' then
              \state\ <= get_wait3796;
            else
              \$1461_lock\ := eclat_true;
              \state\ <= get_pause3797;
            end if;
          when get_wait3805 =>
            if \$1473_lock\(0) = '1' then
              \state\ <= get_wait3805;
            else
              \$1472\ := \$1473\;
              \$v3804\ := \$arr1451_ptr_take\;
              if \$v3804\(0) = '1' then
                \state\ <= q_wait3803;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1472\));
                \state\ <= pause_getI3801;
              end if;
            end if;
          when get_wait3823 =>
            if \$1453_lock\(0) = '1' then
              \state\ <= get_wait3823;
            else
              \$1452\ := \$1453\;
              \$v3822\ := \$arr1451_ptr_take\;
              if \$v3822\(0) = '1' then
                \state\ <= q_wait3821;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1452\));
                \state\ <= pause_getI3819;
              end if;
            end if;
          when get_wait3832 =>
            if \$1459_lock\(0) = '1' then
              \state\ <= get_wait3832;
            else
              \$1458\ := \$1459\;
              \$v3831\ := \$arr1451_ptr_take\;
              if \$v3831\(0) = '1' then
                \state\ <= q_wait3830;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1458\));
                \state\ <= pause_getI3828;
              end if;
            end if;
          when get_wait3837 =>
            if \$1460_lock\(0) = '1' then
              \state\ <= get_wait3837;
            else
              \$1444\ := \$1460\;
              \$v3836\ := \$arr1452_ptr_take\;
              if \$v3836\(0) = '1' then
                \state\ <= q_wait3835;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3833;
              end if;
            end if;
          when get_wait3850 =>
            if \$1481_lock\(0) = '1' then
              \state\ <= get_wait3850;
            else
              \$1480\ := \$1481\;
              \$v3849\ := \$arr1451_ptr_take\;
              if \$v3849\(0) = '1' then
                \state\ <= q_wait3848;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1480\));
                \state\ <= pause_getI3846;
              end if;
            end if;
          when get_wait3859 =>
            if \$1487_lock\(0) = '1' then
              \state\ <= get_wait3859;
            else
              \$1486\ := \$1487\;
              \$v3858\ := \$arr1451_ptr_take\;
              if \$v3858\(0) = '1' then
                \state\ <= q_wait3857;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1486\));
                \state\ <= pause_getI3855;
              end if;
            end if;
          when get_wait3868 =>
            if \$1493_lock\(0) = '1' then
              \state\ <= get_wait3868;
            else
              \$1493_lock\ := eclat_true;
              \state\ <= get_pause3869;
            end if;
          when get_wait3870 =>
            if \$1497_lock\(0) = '1' then
              \state\ <= get_wait3870;
            else
              \$1496\ := \$1497\;
              \$1495\ := \$1496\ & "00000000000000000000000000000001";
              \$1494\ := eclat_sub(\$1495\);
              if \$1493_lock\(0) = '1' then
                \state\ <= get_wait3868;
              else
                \$1493_lock\ := eclat_true;
                \state\ <= get_pause3869;
              end if;
            end if;
          when get_wait3885 =>
            if \$1492_lock\(0) = '1' then
              \state\ <= get_wait3885;
            else
              \$1492_lock\ := eclat_true;
              \state\ <= get_pause3886;
            end if;
          when get_wait3898 =>
            if \$1498_lock\(0) = '1' then
              \state\ <= get_wait3898;
            else
              \$1488_i\ := \$1498\;
              \$v3897\ := eclat_gt(\$1488_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3897\(0) = '1' then
                \$v3896\ := eclat_eq(\$1488_i\ & X"000" & X"15f90");
                if \$v3896\(0) = '1' then
                  \$v3884\ := \$arr1451_ptr_take\;
                  if \$v3884\(0) = '1' then
                    \state\ <= q_wait3883;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3879\ := "00000000000000000000000000000000";
                    \$v3880\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$76_result\ & "0001" & \$v3879\ & "0001" & \$v3880\;
                    \state\ <= pause_setI3881;
                  end if;
                else
                  \$v3895\ := \$arr1451_ptr_take\;
                  if \$v3895\(0) = '1' then
                    \state\ <= q_wait3894;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3891\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$76_result\ & "0010" & \$1488_i\ & "0001" & \$v3891\;
                    \state\ <= pause_setI3892;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811445\;
              end if;
            end if;
          when get_wait3903 =>
            if \$1518_lock\(0) = '1' then
              \state\ <= get_wait3903;
            else
              \$1518_lock\ := eclat_true;
              \state\ <= get_pause3904;
            end if;
          when get_wait3912 =>
            if \$1530_lock\(0) = '1' then
              \state\ <= get_wait3912;
            else
              \$1529\ := \$1530\;
              \$v3911\ := \$arr1451_ptr_take\;
              if \$v3911\(0) = '1' then
                \state\ <= q_wait3910;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1529\));
                \state\ <= pause_getI3908;
              end if;
            end if;
          when get_wait3930 =>
            if \$1510_lock\(0) = '1' then
              \state\ <= get_wait3930;
            else
              \$1509\ := \$1510\;
              \$v3929\ := \$arr1451_ptr_take\;
              if \$v3929\(0) = '1' then
                \state\ <= q_wait3928;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1509\));
                \state\ <= pause_getI3926;
              end if;
            end if;
          when get_wait3939 =>
            if \$1516_lock\(0) = '1' then
              \state\ <= get_wait3939;
            else
              \$1515\ := \$1516\;
              \$v3938\ := \$arr1451_ptr_take\;
              if \$v3938\(0) = '1' then
                \state\ <= q_wait3937;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1515\));
                \state\ <= pause_getI3935;
              end if;
            end if;
          when get_wait3944 =>
            if \$1517_lock\(0) = '1' then
              \state\ <= get_wait3944;
            else
              \$1501\ := \$1517\;
              \$v3943\ := \$arr1452_ptr_take\;
              if \$v3943\(0) = '1' then
                \state\ <= q_wait3942;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3940;
              end if;
            end if;
          when get_wait3957 =>
            if \$1538_lock\(0) = '1' then
              \state\ <= get_wait3957;
            else
              \$1537\ := \$1538\;
              \$v3956\ := \$arr1451_ptr_take\;
              if \$v3956\(0) = '1' then
                \state\ <= q_wait3955;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1537\));
                \state\ <= pause_getI3953;
              end if;
            end if;
          when get_wait3966 =>
            if \$1544_lock\(0) = '1' then
              \state\ <= get_wait3966;
            else
              \$1543\ := \$1544\;
              \$v3965\ := \$arr1451_ptr_take\;
              if \$v3965\(0) = '1' then
                \state\ <= q_wait3964;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1543\));
                \state\ <= pause_getI3962;
              end if;
            end if;
          when get_wait3975 =>
            if \$1550_lock\(0) = '1' then
              \state\ <= get_wait3975;
            else
              \$1550_lock\ := eclat_true;
              \state\ <= get_pause3976;
            end if;
          when get_wait3985 =>
            if \$1549_lock\(0) = '1' then
              \state\ <= get_wait3985;
            else
              \$1549_lock\ := eclat_true;
              \state\ <= get_pause3986;
            end if;
          when get_wait4003 =>
            if \$1551_lock\(0) = '1' then
              \state\ <= get_wait4003;
            else
              \$1545_i\ := \$1551\;
              \$v4002\ := eclat_gt(\$1545_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v4002\(0) = '1' then
                \$v4001\ := eclat_eq(\$1545_i\ & X"000" & X"15f90");
                if \$v4001\(0) = '1' then
                  \$v3984\ := \$arr1451_ptr_take\;
                  if \$v3984\(0) = '1' then
                    \state\ <= q_wait3983;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
                    \state\ <= pause_setI3981;
                  end if;
                else
                  \$v4000\ := \$arr1451_ptr_take\;
                  if \$v4000\(0) = '1' then
                    \state\ <= q_wait3999;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
                    \state\ <= pause_setI3997;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811447\;
              end if;
            end if;
          when get_wait4008 =>
            if \$1571_lock\(0) = '1' then
              \state\ <= get_wait4008;
            else
              \$1571_lock\ := eclat_true;
              \state\ <= get_pause4009;
            end if;
          when get_wait4017 =>
            if \$1583_lock\(0) = '1' then
              \state\ <= get_wait4017;
            else
              \$1582\ := \$1583\;
              \$v4016\ := \$arr1451_ptr_take\;
              if \$v4016\(0) = '1' then
                \state\ <= q_wait4015;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1582\));
                \state\ <= pause_getI4013;
              end if;
            end if;
          when get_wait4035 =>
            if \$1563_lock\(0) = '1' then
              \state\ <= get_wait4035;
            else
              \$1562\ := \$1563\;
              \$v4034\ := \$arr1451_ptr_take\;
              if \$v4034\(0) = '1' then
                \state\ <= q_wait4033;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1562\));
                \state\ <= pause_getI4031;
              end if;
            end if;
          when get_wait4044 =>
            if \$1569_lock\(0) = '1' then
              \state\ <= get_wait4044;
            else
              \$1568\ := \$1569\;
              \$v4043\ := \$arr1451_ptr_take\;
              if \$v4043\(0) = '1' then
                \state\ <= q_wait4042;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1568\));
                \state\ <= pause_getI4040;
              end if;
            end if;
          when get_wait4049 =>
            if \$1570_lock\(0) = '1' then
              \state\ <= get_wait4049;
            else
              \$1554\ := \$1570\;
              \$v4048\ := \$arr1452_ptr_take\;
              if \$v4048\(0) = '1' then
                \state\ <= q_wait4047;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4045;
              end if;
            end if;
          when get_wait4062 =>
            if \$1591_lock\(0) = '1' then
              \state\ <= get_wait4062;
            else
              \$1590\ := \$1591\;
              \$v4061\ := \$arr1451_ptr_take\;
              if \$v4061\(0) = '1' then
                \state\ <= q_wait4060;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1590\));
                \state\ <= pause_getI4058;
              end if;
            end if;
          when get_wait4071 =>
            if \$1597_lock\(0) = '1' then
              \state\ <= get_wait4071;
            else
              \$1596\ := \$1597\;
              \$v4070\ := \$arr1451_ptr_take\;
              if \$v4070\(0) = '1' then
                \state\ <= q_wait4069;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1596\));
                \state\ <= pause_getI4067;
              end if;
            end if;
          when get_wait4076 =>
            if \$1617_lock\(0) = '1' then
              \state\ <= get_wait4076;
            else
              \$1617_lock\ := eclat_true;
              \state\ <= get_pause4077;
            end if;
          when get_wait4085 =>
            if \$1629_lock\(0) = '1' then
              \state\ <= get_wait4085;
            else
              \$1628\ := \$1629\;
              \$v4084\ := \$arr1451_ptr_take\;
              if \$v4084\(0) = '1' then
                \state\ <= q_wait4083;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1628\));
                \state\ <= pause_getI4081;
              end if;
            end if;
          when get_wait4103 =>
            if \$1609_lock\(0) = '1' then
              \state\ <= get_wait4103;
            else
              \$1608\ := \$1609\;
              \$v4102\ := \$arr1451_ptr_take\;
              if \$v4102\(0) = '1' then
                \state\ <= q_wait4101;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1608\));
                \state\ <= pause_getI4099;
              end if;
            end if;
          when get_wait4112 =>
            if \$1615_lock\(0) = '1' then
              \state\ <= get_wait4112;
            else
              \$1614\ := \$1615\;
              \$v4111\ := \$arr1451_ptr_take\;
              if \$v4111\(0) = '1' then
                \state\ <= q_wait4110;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1614\));
                \state\ <= pause_getI4108;
              end if;
            end if;
          when get_wait4117 =>
            if \$1616_lock\(0) = '1' then
              \state\ <= get_wait4117;
            else
              \$1600\ := \$1616\;
              \$v4116\ := \$arr1452_ptr_take\;
              if \$v4116\(0) = '1' then
                \state\ <= q_wait4115;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4113;
              end if;
            end if;
          when get_wait4130 =>
            if \$1637_lock\(0) = '1' then
              \state\ <= get_wait4130;
            else
              \$1636\ := \$1637\;
              \$v4129\ := \$arr1451_ptr_take\;
              if \$v4129\(0) = '1' then
                \state\ <= q_wait4128;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1636\));
                \state\ <= pause_getI4126;
              end if;
            end if;
          when get_wait4139 =>
            if \$1643_lock\(0) = '1' then
              \state\ <= get_wait4139;
            else
              \$1642\ := \$1643\;
              \$v4138\ := \$arr1451_ptr_take\;
              if \$v4138\(0) = '1' then
                \state\ <= q_wait4137;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1642\));
                \state\ <= pause_getI4135;
              end if;
            end if;
          when get_wait4144 =>
            if \$1663_lock\(0) = '1' then
              \state\ <= get_wait4144;
            else
              \$1663_lock\ := eclat_true;
              \state\ <= get_pause4145;
            end if;
          when get_wait4153 =>
            if \$1675_lock\(0) = '1' then
              \state\ <= get_wait4153;
            else
              \$1674\ := \$1675\;
              \$v4152\ := \$arr1451_ptr_take\;
              if \$v4152\(0) = '1' then
                \state\ <= q_wait4151;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1674\));
                \state\ <= pause_getI4149;
              end if;
            end if;
          when get_wait4171 =>
            if \$1655_lock\(0) = '1' then
              \state\ <= get_wait4171;
            else
              \$1654\ := \$1655\;
              \$v4170\ := \$arr1451_ptr_take\;
              if \$v4170\(0) = '1' then
                \state\ <= q_wait4169;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1654\));
                \state\ <= pause_getI4167;
              end if;
            end if;
          when get_wait4180 =>
            if \$1661_lock\(0) = '1' then
              \state\ <= get_wait4180;
            else
              \$1660\ := \$1661\;
              \$v4179\ := \$arr1451_ptr_take\;
              if \$v4179\(0) = '1' then
                \state\ <= q_wait4178;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1660\));
                \state\ <= pause_getI4176;
              end if;
            end if;
          when get_wait4185 =>
            if \$1662_lock\(0) = '1' then
              \state\ <= get_wait4185;
            else
              \$1646\ := \$1662\;
              \$v4184\ := \$arr1452_ptr_take\;
              if \$v4184\(0) = '1' then
                \state\ <= q_wait4183;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4181;
              end if;
            end if;
          when get_wait4198 =>
            if \$1683_lock\(0) = '1' then
              \state\ <= get_wait4198;
            else
              \$1682\ := \$1683\;
              \$v4197\ := \$arr1451_ptr_take\;
              if \$v4197\(0) = '1' then
                \state\ <= q_wait4196;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1682\));
                \state\ <= pause_getI4194;
              end if;
            end if;
          when get_wait4207 =>
            if \$1689_lock\(0) = '1' then
              \state\ <= get_wait4207;
            else
              \$1688\ := \$1689\;
              \$v4206\ := \$arr1451_ptr_take\;
              if \$v4206\(0) = '1' then
                \state\ <= q_wait4205;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1688\));
                \state\ <= pause_getI4203;
              end if;
            end if;
          when get_wait4216 =>
            if \$v16_lock\(0) = '1' then
              \state\ <= get_wait4216;
            else
              \$v17\ := \$v16\;
              \$v4215\ := \$arr1451_ptr_take\;
              if \$v4215\(0) = '1' then
                \state\ <= q_wait4214;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v17\));
                \state\ <= pause_getI4212;
              end if;
            end if;
          when pause_getI1464 =>
            \state\ <= pause_getII1465;
          when pause_getI1468 =>
            \state\ <= pause_getII1469;
          when pause_getI1480 =>
            \state\ <= pause_getII1481;
          when pause_getI1492 =>
            \state\ <= pause_getII1493;
          when pause_getI1508 =>
            \state\ <= pause_getII1509;
          when pause_getI1513 =>
            \state\ <= pause_getII1514;
          when pause_getI1517 =>
            \state\ <= pause_getII1518;
          when pause_getI1526 =>
            \state\ <= pause_getII1527;
          when pause_getI1531 =>
            \state\ <= pause_getII1532;
          when pause_getI1535 =>
            \state\ <= pause_getII1536;
          when pause_getI1540 =>
            \state\ <= pause_getII1541;
          when pause_getI1545 =>
            \state\ <= pause_getII1546;
          when pause_getI1553 =>
            \state\ <= pause_getII1554;
          when pause_getI1558 =>
            \state\ <= pause_getII1559;
          when pause_getI1562 =>
            \state\ <= pause_getII1563;
          when pause_getI1567 =>
            \state\ <= pause_getII1568;
          when pause_getI1576 =>
            \state\ <= pause_getII1577;
          when pause_getI1581 =>
            \state\ <= pause_getII1582;
          when pause_getI1585 =>
            \state\ <= pause_getII1586;
          when pause_getI1594 =>
            \state\ <= pause_getII1595;
          when pause_getI1599 =>
            \state\ <= pause_getII1600;
          when pause_getI1603 =>
            \state\ <= pause_getII1604;
          when pause_getI1608 =>
            \state\ <= pause_getII1609;
          when pause_getI1613 =>
            \state\ <= pause_getII1614;
          when pause_getI1621 =>
            \state\ <= pause_getII1622;
          when pause_getI1626 =>
            \state\ <= pause_getII1627;
          when pause_getI1630 =>
            \state\ <= pause_getII1631;
          when pause_getI1635 =>
            \state\ <= pause_getII1636;
          when pause_getI1646 =>
            \state\ <= pause_getII1647;
          when pause_getI1650 =>
            \state\ <= pause_getII1651;
          when pause_getI1662 =>
            \state\ <= pause_getII1663;
          when pause_getI1674 =>
            \state\ <= pause_getII1675;
          when pause_getI1690 =>
            \state\ <= pause_getII1691;
          when pause_getI1695 =>
            \state\ <= pause_getII1696;
          when pause_getI1699 =>
            \state\ <= pause_getII1700;
          when pause_getI1708 =>
            \state\ <= pause_getII1709;
          when pause_getI1713 =>
            \state\ <= pause_getII1714;
          when pause_getI1717 =>
            \state\ <= pause_getII1718;
          when pause_getI1722 =>
            \state\ <= pause_getII1723;
          when pause_getI1727 =>
            \state\ <= pause_getII1728;
          when pause_getI1735 =>
            \state\ <= pause_getII1736;
          when pause_getI1740 =>
            \state\ <= pause_getII1741;
          when pause_getI1744 =>
            \state\ <= pause_getII1745;
          when pause_getI1749 =>
            \state\ <= pause_getII1750;
          when pause_getI1758 =>
            \state\ <= pause_getII1759;
          when pause_getI1763 =>
            \state\ <= pause_getII1764;
          when pause_getI1767 =>
            \state\ <= pause_getII1768;
          when pause_getI1776 =>
            \state\ <= pause_getII1777;
          when pause_getI1781 =>
            \state\ <= pause_getII1782;
          when pause_getI1785 =>
            \state\ <= pause_getII1786;
          when pause_getI1790 =>
            \state\ <= pause_getII1791;
          when pause_getI1795 =>
            \state\ <= pause_getII1796;
          when pause_getI1803 =>
            \state\ <= pause_getII1804;
          when pause_getI1808 =>
            \state\ <= pause_getII1809;
          when pause_getI1812 =>
            \state\ <= pause_getII1813;
          when pause_getI1817 =>
            \state\ <= pause_getII1818;
          when pause_getI1828 =>
            \state\ <= pause_getII1829;
          when pause_getI1832 =>
            \state\ <= pause_getII1833;
          when pause_getI1844 =>
            \state\ <= pause_getII1845;
          when pause_getI1856 =>
            \state\ <= pause_getII1857;
          when pause_getI1872 =>
            \state\ <= pause_getII1873;
          when pause_getI1877 =>
            \state\ <= pause_getII1878;
          when pause_getI1881 =>
            \state\ <= pause_getII1882;
          when pause_getI1890 =>
            \state\ <= pause_getII1891;
          when pause_getI1895 =>
            \state\ <= pause_getII1896;
          when pause_getI1899 =>
            \state\ <= pause_getII1900;
          when pause_getI1904 =>
            \state\ <= pause_getII1905;
          when pause_getI1909 =>
            \state\ <= pause_getII1910;
          when pause_getI1917 =>
            \state\ <= pause_getII1918;
          when pause_getI1922 =>
            \state\ <= pause_getII1923;
          when pause_getI1926 =>
            \state\ <= pause_getII1927;
          when pause_getI1931 =>
            \state\ <= pause_getII1932;
          when pause_getI1940 =>
            \state\ <= pause_getII1941;
          when pause_getI1945 =>
            \state\ <= pause_getII1946;
          when pause_getI1949 =>
            \state\ <= pause_getII1950;
          when pause_getI1958 =>
            \state\ <= pause_getII1959;
          when pause_getI1963 =>
            \state\ <= pause_getII1964;
          when pause_getI1967 =>
            \state\ <= pause_getII1968;
          when pause_getI1972 =>
            \state\ <= pause_getII1973;
          when pause_getI1977 =>
            \state\ <= pause_getII1978;
          when pause_getI1985 =>
            \state\ <= pause_getII1986;
          when pause_getI1990 =>
            \state\ <= pause_getII1991;
          when pause_getI1994 =>
            \state\ <= pause_getII1995;
          when pause_getI1999 =>
            \state\ <= pause_getII2000;
          when pause_getI2010 =>
            \state\ <= pause_getII2011;
          when pause_getI2014 =>
            \state\ <= pause_getII2015;
          when pause_getI2026 =>
            \state\ <= pause_getII2027;
          when pause_getI2038 =>
            \state\ <= pause_getII2039;
          when pause_getI2054 =>
            \state\ <= pause_getII2055;
          when pause_getI2059 =>
            \state\ <= pause_getII2060;
          when pause_getI2063 =>
            \state\ <= pause_getII2064;
          when pause_getI2072 =>
            \state\ <= pause_getII2073;
          when pause_getI2077 =>
            \state\ <= pause_getII2078;
          when pause_getI2081 =>
            \state\ <= pause_getII2082;
          when pause_getI2086 =>
            \state\ <= pause_getII2087;
          when pause_getI2091 =>
            \state\ <= pause_getII2092;
          when pause_getI2099 =>
            \state\ <= pause_getII2100;
          when pause_getI2104 =>
            \state\ <= pause_getII2105;
          when pause_getI2108 =>
            \state\ <= pause_getII2109;
          when pause_getI2113 =>
            \state\ <= pause_getII2114;
          when pause_getI2122 =>
            \state\ <= pause_getII2123;
          when pause_getI2127 =>
            \state\ <= pause_getII2128;
          when pause_getI2131 =>
            \state\ <= pause_getII2132;
          when pause_getI2140 =>
            \state\ <= pause_getII2141;
          when pause_getI2145 =>
            \state\ <= pause_getII2146;
          when pause_getI2149 =>
            \state\ <= pause_getII2150;
          when pause_getI2154 =>
            \state\ <= pause_getII2155;
          when pause_getI2159 =>
            \state\ <= pause_getII2160;
          when pause_getI2167 =>
            \state\ <= pause_getII2168;
          when pause_getI2172 =>
            \state\ <= pause_getII2173;
          when pause_getI2176 =>
            \state\ <= pause_getII2177;
          when pause_getI2181 =>
            \state\ <= pause_getII2182;
          when pause_getI2191 =>
            \state\ <= pause_getII2192;
          when pause_getI2207 =>
            \state\ <= pause_getII2208;
          when pause_getI2230 =>
            \state\ <= pause_getII2231;
          when pause_getI2245 =>
            \state\ <= pause_getII2246;
          when pause_getI2250 =>
            \state\ <= pause_getII2251;
          when pause_getI2254 =>
            \state\ <= pause_getII2255;
          when pause_getI2263 =>
            \state\ <= pause_getII2264;
          when pause_getI2268 =>
            \state\ <= pause_getII2269;
          when pause_getI2272 =>
            \state\ <= pause_getII2273;
          when pause_getI2277 =>
            \state\ <= pause_getII2278;
          when pause_getI2282 =>
            \state\ <= pause_getII2283;
          when pause_getI2290 =>
            \state\ <= pause_getII2291;
          when pause_getI2295 =>
            \state\ <= pause_getII2296;
          when pause_getI2299 =>
            \state\ <= pause_getII2300;
          when pause_getI2304 =>
            \state\ <= pause_getII2305;
          when pause_getI2313 =>
            \state\ <= pause_getII2314;
          when pause_getI2318 =>
            \state\ <= pause_getII2319;
          when pause_getI2322 =>
            \state\ <= pause_getII2323;
          when pause_getI2331 =>
            \state\ <= pause_getII2332;
          when pause_getI2336 =>
            \state\ <= pause_getII2337;
          when pause_getI2340 =>
            \state\ <= pause_getII2341;
          when pause_getI2345 =>
            \state\ <= pause_getII2346;
          when pause_getI2350 =>
            \state\ <= pause_getII2351;
          when pause_getI2358 =>
            \state\ <= pause_getII2359;
          when pause_getI2363 =>
            \state\ <= pause_getII2364;
          when pause_getI2367 =>
            \state\ <= pause_getII2368;
          when pause_getI2372 =>
            \state\ <= pause_getII2373;
          when pause_getI2382 =>
            \state\ <= pause_getII2383;
          when pause_getI2398 =>
            \state\ <= pause_getII2399;
          when pause_getI2421 =>
            \state\ <= pause_getII2422;
          when pause_getI2439 =>
            \state\ <= pause_getII2440;
          when pause_getI2444 =>
            \state\ <= pause_getII2445;
          when pause_getI2448 =>
            \state\ <= pause_getII2449;
          when pause_getI2457 =>
            \state\ <= pause_getII2458;
          when pause_getI2462 =>
            \state\ <= pause_getII2463;
          when pause_getI2466 =>
            \state\ <= pause_getII2467;
          when pause_getI2471 =>
            \state\ <= pause_getII2472;
          when pause_getI2476 =>
            \state\ <= pause_getII2477;
          when pause_getI2484 =>
            \state\ <= pause_getII2485;
          when pause_getI2489 =>
            \state\ <= pause_getII2490;
          when pause_getI2493 =>
            \state\ <= pause_getII2494;
          when pause_getI2498 =>
            \state\ <= pause_getII2499;
          when pause_getI2507 =>
            \state\ <= pause_getII2508;
          when pause_getI2512 =>
            \state\ <= pause_getII2513;
          when pause_getI2516 =>
            \state\ <= pause_getII2517;
          when pause_getI2525 =>
            \state\ <= pause_getII2526;
          when pause_getI2530 =>
            \state\ <= pause_getII2531;
          when pause_getI2534 =>
            \state\ <= pause_getII2535;
          when pause_getI2539 =>
            \state\ <= pause_getII2540;
          when pause_getI2544 =>
            \state\ <= pause_getII2545;
          when pause_getI2552 =>
            \state\ <= pause_getII2553;
          when pause_getI2557 =>
            \state\ <= pause_getII2558;
          when pause_getI2561 =>
            \state\ <= pause_getII2562;
          when pause_getI2566 =>
            \state\ <= pause_getII2567;
          when pause_getI2576 =>
            \state\ <= pause_getII2577;
          when pause_getI2586 =>
            \state\ <= pause_getII2587;
          when pause_getI2603 =>
            \state\ <= pause_getII2604;
          when pause_getI2608 =>
            \state\ <= pause_getII2609;
          when pause_getI2619 =>
            \state\ <= pause_getII2620;
          when pause_getI2624 =>
            \state\ <= pause_getII2625;
          when pause_getI2628 =>
            \state\ <= pause_getII2629;
          when pause_getI2637 =>
            \state\ <= pause_getII2638;
          when pause_getI2642 =>
            \state\ <= pause_getII2643;
          when pause_getI2646 =>
            \state\ <= pause_getII2647;
          when pause_getI2651 =>
            \state\ <= pause_getII2652;
          when pause_getI2656 =>
            \state\ <= pause_getII2657;
          when pause_getI2664 =>
            \state\ <= pause_getII2665;
          when pause_getI2669 =>
            \state\ <= pause_getII2670;
          when pause_getI2673 =>
            \state\ <= pause_getII2674;
          when pause_getI2678 =>
            \state\ <= pause_getII2679;
          when pause_getI2687 =>
            \state\ <= pause_getII2688;
          when pause_getI2692 =>
            \state\ <= pause_getII2693;
          when pause_getI2696 =>
            \state\ <= pause_getII2697;
          when pause_getI2705 =>
            \state\ <= pause_getII2706;
          when pause_getI2710 =>
            \state\ <= pause_getII2711;
          when pause_getI2714 =>
            \state\ <= pause_getII2715;
          when pause_getI2719 =>
            \state\ <= pause_getII2720;
          when pause_getI2724 =>
            \state\ <= pause_getII2725;
          when pause_getI2732 =>
            \state\ <= pause_getII2733;
          when pause_getI2737 =>
            \state\ <= pause_getII2738;
          when pause_getI2741 =>
            \state\ <= pause_getII2742;
          when pause_getI2746 =>
            \state\ <= pause_getII2747;
          when pause_getI2756 =>
            \state\ <= pause_getII2757;
          when pause_getI2766 =>
            \state\ <= pause_getII2767;
          when pause_getI2783 =>
            \state\ <= pause_getII2784;
          when pause_getI2788 =>
            \state\ <= pause_getII2789;
          when pause_getI2799 =>
            \state\ <= pause_getII2800;
          when pause_getI2804 =>
            \state\ <= pause_getII2805;
          when pause_getI2808 =>
            \state\ <= pause_getII2809;
          when pause_getI2817 =>
            \state\ <= pause_getII2818;
          when pause_getI2822 =>
            \state\ <= pause_getII2823;
          when pause_getI2826 =>
            \state\ <= pause_getII2827;
          when pause_getI2831 =>
            \state\ <= pause_getII2832;
          when pause_getI2836 =>
            \state\ <= pause_getII2837;
          when pause_getI2844 =>
            \state\ <= pause_getII2845;
          when pause_getI2849 =>
            \state\ <= pause_getII2850;
          when pause_getI2853 =>
            \state\ <= pause_getII2854;
          when pause_getI2858 =>
            \state\ <= pause_getII2859;
          when pause_getI2867 =>
            \state\ <= pause_getII2868;
          when pause_getI2872 =>
            \state\ <= pause_getII2873;
          when pause_getI2876 =>
            \state\ <= pause_getII2877;
          when pause_getI2885 =>
            \state\ <= pause_getII2886;
          when pause_getI2890 =>
            \state\ <= pause_getII2891;
          when pause_getI2894 =>
            \state\ <= pause_getII2895;
          when pause_getI2899 =>
            \state\ <= pause_getII2900;
          when pause_getI2904 =>
            \state\ <= pause_getII2905;
          when pause_getI2912 =>
            \state\ <= pause_getII2913;
          when pause_getI2917 =>
            \state\ <= pause_getII2918;
          when pause_getI2921 =>
            \state\ <= pause_getII2922;
          when pause_getI2926 =>
            \state\ <= pause_getII2927;
          when pause_getI2936 =>
            \state\ <= pause_getII2937;
          when pause_getI2946 =>
            \state\ <= pause_getII2947;
          when pause_getI2963 =>
            \state\ <= pause_getII2964;
          when pause_getI2968 =>
            \state\ <= pause_getII2969;
          when pause_getI2979 =>
            \state\ <= pause_getII2980;
          when pause_getI2984 =>
            \state\ <= pause_getII2985;
          when pause_getI2988 =>
            \state\ <= pause_getII2989;
          when pause_getI2997 =>
            \state\ <= pause_getII2998;
          when pause_getI3002 =>
            \state\ <= pause_getII3003;
          when pause_getI3006 =>
            \state\ <= pause_getII3007;
          when pause_getI3011 =>
            \state\ <= pause_getII3012;
          when pause_getI3016 =>
            \state\ <= pause_getII3017;
          when pause_getI3024 =>
            \state\ <= pause_getII3025;
          when pause_getI3029 =>
            \state\ <= pause_getII3030;
          when pause_getI3033 =>
            \state\ <= pause_getII3034;
          when pause_getI3038 =>
            \state\ <= pause_getII3039;
          when pause_getI3047 =>
            \state\ <= pause_getII3048;
          when pause_getI3052 =>
            \state\ <= pause_getII3053;
          when pause_getI3056 =>
            \state\ <= pause_getII3057;
          when pause_getI3065 =>
            \state\ <= pause_getII3066;
          when pause_getI3070 =>
            \state\ <= pause_getII3071;
          when pause_getI3074 =>
            \state\ <= pause_getII3075;
          when pause_getI3079 =>
            \state\ <= pause_getII3080;
          when pause_getI3084 =>
            \state\ <= pause_getII3085;
          when pause_getI3092 =>
            \state\ <= pause_getII3093;
          when pause_getI3097 =>
            \state\ <= pause_getII3098;
          when pause_getI3101 =>
            \state\ <= pause_getII3102;
          when pause_getI3106 =>
            \state\ <= pause_getII3107;
          when pause_getI3117 =>
            \state\ <= pause_getII3118;
          when pause_getI3121 =>
            \state\ <= pause_getII3122;
          when pause_getI3133 =>
            \state\ <= pause_getII3134;
          when pause_getI3145 =>
            \state\ <= pause_getII3146;
          when pause_getI3150 =>
            \state\ <= pause_getII3151;
          when pause_getI3161 =>
            \state\ <= pause_getII3162;
          when pause_getI3166 =>
            \state\ <= pause_getII3167;
          when pause_getI3170 =>
            \state\ <= pause_getII3171;
          when pause_getI3179 =>
            \state\ <= pause_getII3180;
          when pause_getI3184 =>
            \state\ <= pause_getII3185;
          when pause_getI3188 =>
            \state\ <= pause_getII3189;
          when pause_getI3193 =>
            \state\ <= pause_getII3194;
          when pause_getI3198 =>
            \state\ <= pause_getII3199;
          when pause_getI3206 =>
            \state\ <= pause_getII3207;
          when pause_getI3211 =>
            \state\ <= pause_getII3212;
          when pause_getI3215 =>
            \state\ <= pause_getII3216;
          when pause_getI3220 =>
            \state\ <= pause_getII3221;
          when pause_getI3231 =>
            \state\ <= pause_getII3232;
          when pause_getI3235 =>
            \state\ <= pause_getII3236;
          when pause_getI3247 =>
            \state\ <= pause_getII3248;
          when pause_getI3259 =>
            \state\ <= pause_getII3260;
          when pause_getI3264 =>
            \state\ <= pause_getII3265;
          when pause_getI3275 =>
            \state\ <= pause_getII3276;
          when pause_getI3280 =>
            \state\ <= pause_getII3281;
          when pause_getI3284 =>
            \state\ <= pause_getII3285;
          when pause_getI3293 =>
            \state\ <= pause_getII3294;
          when pause_getI3298 =>
            \state\ <= pause_getII3299;
          when pause_getI3302 =>
            \state\ <= pause_getII3303;
          when pause_getI3307 =>
            \state\ <= pause_getII3308;
          when pause_getI3312 =>
            \state\ <= pause_getII3313;
          when pause_getI3320 =>
            \state\ <= pause_getII3321;
          when pause_getI3325 =>
            \state\ <= pause_getII3326;
          when pause_getI3329 =>
            \state\ <= pause_getII3330;
          when pause_getI3334 =>
            \state\ <= pause_getII3335;
          when pause_getI3345 =>
            \state\ <= pause_getII3346;
          when pause_getI3349 =>
            \state\ <= pause_getII3350;
          when pause_getI3361 =>
            \state\ <= pause_getII3362;
          when pause_getI3373 =>
            \state\ <= pause_getII3374;
          when pause_getI3378 =>
            \state\ <= pause_getII3379;
          when pause_getI3389 =>
            \state\ <= pause_getII3390;
          when pause_getI3394 =>
            \state\ <= pause_getII3395;
          when pause_getI3398 =>
            \state\ <= pause_getII3399;
          when pause_getI3407 =>
            \state\ <= pause_getII3408;
          when pause_getI3412 =>
            \state\ <= pause_getII3413;
          when pause_getI3416 =>
            \state\ <= pause_getII3417;
          when pause_getI3421 =>
            \state\ <= pause_getII3422;
          when pause_getI3426 =>
            \state\ <= pause_getII3427;
          when pause_getI3434 =>
            \state\ <= pause_getII3435;
          when pause_getI3439 =>
            \state\ <= pause_getII3440;
          when pause_getI3443 =>
            \state\ <= pause_getII3444;
          when pause_getI3448 =>
            \state\ <= pause_getII3449;
          when pause_getI3458 =>
            \state\ <= pause_getII3459;
          when pause_getI3468 =>
            \state\ <= pause_getII3469;
          when pause_getI3485 =>
            \state\ <= pause_getII3486;
          when pause_getI3503 =>
            \state\ <= pause_getII3504;
          when pause_getI3508 =>
            \state\ <= pause_getII3509;
          when pause_getI3512 =>
            \state\ <= pause_getII3513;
          when pause_getI3521 =>
            \state\ <= pause_getII3522;
          when pause_getI3526 =>
            \state\ <= pause_getII3527;
          when pause_getI3530 =>
            \state\ <= pause_getII3531;
          when pause_getI3535 =>
            \state\ <= pause_getII3536;
          when pause_getI3540 =>
            \state\ <= pause_getII3541;
          when pause_getI3548 =>
            \state\ <= pause_getII3549;
          when pause_getI3553 =>
            \state\ <= pause_getII3554;
          when pause_getI3557 =>
            \state\ <= pause_getII3558;
          when pause_getI3562 =>
            \state\ <= pause_getII3563;
          when pause_getI3572 =>
            \state\ <= pause_getII3573;
          when pause_getI3583 =>
            \state\ <= pause_getII3584;
          when pause_getI3601 =>
            \state\ <= pause_getII3602;
          when pause_getI3605 =>
            \state\ <= pause_getII3606;
          when pause_getI3610 =>
            \state\ <= pause_getII3611;
          when pause_getI3615 =>
            \state\ <= pause_getII3616;
          when pause_getI3626 =>
            \state\ <= pause_getII3627;
          when pause_getI3631 =>
            \state\ <= pause_getII3632;
          when pause_getI3635 =>
            \state\ <= pause_getII3636;
          when pause_getI3644 =>
            \state\ <= pause_getII3645;
          when pause_getI3649 =>
            \state\ <= pause_getII3650;
          when pause_getI3653 =>
            \state\ <= pause_getII3654;
          when pause_getI3658 =>
            \state\ <= pause_getII3659;
          when pause_getI3663 =>
            \state\ <= pause_getII3664;
          when pause_getI3671 =>
            \state\ <= pause_getII3672;
          when pause_getI3676 =>
            \state\ <= pause_getII3677;
          when pause_getI3680 =>
            \state\ <= pause_getII3681;
          when pause_getI3685 =>
            \state\ <= pause_getII3686;
          when pause_getI3696 =>
            \state\ <= pause_getII3697;
          when pause_getI3700 =>
            \state\ <= pause_getII3701;
          when pause_getI3712 =>
            \state\ <= pause_getII3713;
          when pause_getI3724 =>
            \state\ <= pause_getII3725;
          when pause_getI3733 =>
            \state\ <= pause_getII3734;
          when pause_getI3738 =>
            \state\ <= pause_getII3739;
          when pause_getI3742 =>
            \state\ <= pause_getII3743;
          when pause_getI3751 =>
            \state\ <= pause_getII3752;
          when pause_getI3756 =>
            \state\ <= pause_getII3757;
          when pause_getI3760 =>
            \state\ <= pause_getII3761;
          when pause_getI3765 =>
            \state\ <= pause_getII3766;
          when pause_getI3770 =>
            \state\ <= pause_getII3771;
          when pause_getI3778 =>
            \state\ <= pause_getII3779;
          when pause_getI3783 =>
            \state\ <= pause_getII3784;
          when pause_getI3787 =>
            \state\ <= pause_getII3788;
          when pause_getI3792 =>
            \state\ <= pause_getII3793;
          when pause_getI3801 =>
            \state\ <= pause_getII3802;
          when pause_getI3806 =>
            \state\ <= pause_getII3807;
          when pause_getI3810 =>
            \state\ <= pause_getII3811;
          when pause_getI3819 =>
            \state\ <= pause_getII3820;
          when pause_getI3824 =>
            \state\ <= pause_getII3825;
          when pause_getI3828 =>
            \state\ <= pause_getII3829;
          when pause_getI3833 =>
            \state\ <= pause_getII3834;
          when pause_getI3838 =>
            \state\ <= pause_getII3839;
          when pause_getI3846 =>
            \state\ <= pause_getII3847;
          when pause_getI3851 =>
            \state\ <= pause_getII3852;
          when pause_getI3855 =>
            \state\ <= pause_getII3856;
          when pause_getI3860 =>
            \state\ <= pause_getII3861;
          when pause_getI3871 =>
            \state\ <= pause_getII3872;
          when pause_getI3875 =>
            \state\ <= pause_getII3876;
          when pause_getI3887 =>
            \state\ <= pause_getII3888;
          when pause_getI3899 =>
            \state\ <= pause_getII3900;
          when pause_getI3908 =>
            \state\ <= pause_getII3909;
          when pause_getI3913 =>
            \state\ <= pause_getII3914;
          when pause_getI3917 =>
            \state\ <= pause_getII3918;
          when pause_getI3926 =>
            \state\ <= pause_getII3927;
          when pause_getI3931 =>
            \state\ <= pause_getII3932;
          when pause_getI3935 =>
            \state\ <= pause_getII3936;
          when pause_getI3940 =>
            \state\ <= pause_getII3941;
          when pause_getI3945 =>
            \state\ <= pause_getII3946;
          when pause_getI3953 =>
            \state\ <= pause_getII3954;
          when pause_getI3958 =>
            \state\ <= pause_getII3959;
          when pause_getI3962 =>
            \state\ <= pause_getII3963;
          when pause_getI3967 =>
            \state\ <= pause_getII3968;
          when pause_getI3977 =>
            \state\ <= pause_getII3978;
          when pause_getI3987 =>
            \state\ <= pause_getII3988;
          when pause_getI4004 =>
            \state\ <= pause_getII4005;
          when pause_getI4013 =>
            \state\ <= pause_getII4014;
          when pause_getI4018 =>
            \state\ <= pause_getII4019;
          when pause_getI4022 =>
            \state\ <= pause_getII4023;
          when pause_getI4031 =>
            \state\ <= pause_getII4032;
          when pause_getI4036 =>
            \state\ <= pause_getII4037;
          when pause_getI4040 =>
            \state\ <= pause_getII4041;
          when pause_getI4045 =>
            \state\ <= pause_getII4046;
          when pause_getI4050 =>
            \state\ <= pause_getII4051;
          when pause_getI4058 =>
            \state\ <= pause_getII4059;
          when pause_getI4063 =>
            \state\ <= pause_getII4064;
          when pause_getI4067 =>
            \state\ <= pause_getII4068;
          when pause_getI4072 =>
            \state\ <= pause_getII4073;
          when pause_getI4081 =>
            \state\ <= pause_getII4082;
          when pause_getI4086 =>
            \state\ <= pause_getII4087;
          when pause_getI4090 =>
            \state\ <= pause_getII4091;
          when pause_getI4099 =>
            \state\ <= pause_getII4100;
          when pause_getI4104 =>
            \state\ <= pause_getII4105;
          when pause_getI4108 =>
            \state\ <= pause_getII4109;
          when pause_getI4113 =>
            \state\ <= pause_getII4114;
          when pause_getI4118 =>
            \state\ <= pause_getII4119;
          when pause_getI4126 =>
            \state\ <= pause_getII4127;
          when pause_getI4131 =>
            \state\ <= pause_getII4132;
          when pause_getI4135 =>
            \state\ <= pause_getII4136;
          when pause_getI4140 =>
            \state\ <= pause_getII4141;
          when pause_getI4149 =>
            \state\ <= pause_getII4150;
          when pause_getI4154 =>
            \state\ <= pause_getII4155;
          when pause_getI4158 =>
            \state\ <= pause_getII4159;
          when pause_getI4167 =>
            \state\ <= pause_getII4168;
          when pause_getI4172 =>
            \state\ <= pause_getII4173;
          when pause_getI4176 =>
            \state\ <= pause_getII4177;
          when pause_getI4181 =>
            \state\ <= pause_getII4182;
          when pause_getI4186 =>
            \state\ <= pause_getII4187;
          when pause_getI4194 =>
            \state\ <= pause_getII4195;
          when pause_getI4199 =>
            \state\ <= pause_getII4200;
          when pause_getI4203 =>
            \state\ <= pause_getII4204;
          when pause_getI4208 =>
            \state\ <= pause_getII4209;
          when pause_getI4212 =>
            \state\ <= pause_getII4213;
          when pause_getI4217 =>
            \state\ <= pause_getII4218;
          when pause_getII1465 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v73\ := \$arr1452_value\;
            if \$v73_lock\(0) = '1' then
              \state\ <= get_wait1463;
            else
              \$v74\ := \$v73\;
              \$v75\ := \$v74\ & "00000000000000000000000000000001";
              \$v77\ := eclat_sub(\$v75\);
              if \$v76_lock\(0) = '1' then
                \state\ <= get_wait1461;
              else
                \$v76_lock\ := eclat_true;
                \state\ <= get_pause1462;
              end if;
            end if;
          when pause_getII1469 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1467\ := \$arr1452_ptr_take\;
            if \$v1467\(0) = '1' then
              \state\ <= q_wait1466;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1464;
            end if;
          when pause_getII1481 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$v67_lock\(0) = '1' then
              \state\ <= get_wait1478;
            else
              \$v67_lock\ := eclat_true;
              \state\ <= get_pause1479;
            end if;
          when pause_getII1493 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v60\ := \$arr1452_value\;
            if \$v60_lock\(0) = '1' then
              \state\ <= get_wait1491;
            else
              \$81_i\ := \$v60\;
              \$v1490\ := eclat_gt(\$81_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1490\(0) = '1' then
                \$v1489\ := eclat_eq(\$81_i\ & X"000" & X"15f90");
                if \$v1489\(0) = '1' then
                  \$v1477\ := \$arr1451_ptr_take\;
                  if \$v1477\(0) = '1' then
                    \state\ <= q_wait1476;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1472\ := "00000000000000000000000000000000";
                    \$v1473\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$71_result_after_f\ & "0001" & \$v1472\ & "0001" & \$v1473\;
                    \state\ <= pause_setI1474;
                  end if;
                else
                  \$v1488\ := \$arr1451_ptr_take\;
                  if \$v1488\(0) = '1' then
                    \state\ <= q_wait1487;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1484\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$71_result_after_f\ & "0010" & \$81_i\ & "0001" & \$v1484\;
                    \state\ <= pause_setI1485;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811388\;
              end if;
            end if;
          when pause_getII1509 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v41\ := \$arr1451_value\;
            \$v42\ := \$v41\(36 to 71);
            \$v1506\ := \$v42\;
            \$v1507\ := \$v1506\(0 to 3);
            \$v1505\ := \$v1506\(4 to 35);
            case \$v1507\ is
            when "0010" =>
              \$137_i\ := \$v1505\(0 to 31);
              \$v44\ := \$137_i\;
              if \$v43_lock\(0) = '1' then
                \state\ <= get_wait1503;
              else
                \$v43_lock\ := eclat_true;
                \state\ <= get_pause1504;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811391\;
            end case;
          when pause_getII1514 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v39\ := \$arr1452_value\;
            if \$v39_lock\(0) = '1' then
              \state\ <= get_wait1512;
            else
              \$v40\ := \$v39\;
              \$v1511\ := \$arr1451_ptr_take\;
              if \$v1511\(0) = '1' then
                \state\ <= q_wait1510;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v40\));
                \state\ <= pause_getI1508;
              end if;
            end if;
          when pause_getII1518 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1516\ := \$arr1452_ptr_take\;
            if \$v1516\(0) = '1' then
              \state\ <= q_wait1515;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1513;
            end if;
          when pause_getII1527 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v33\ := \$arr1451_value\;
            \$v36\ := \$v33\(72 to 107);
            \$v1525\ := "00000000000000000000000000000000";
            \$v38\ := "0000" & \$v1525\ & \$v35\ & \$v36\;
            \$v1524\ := \$arr1451_ptr_take\;
            if \$v1524\(0) = '1' then
              \state\ <= q_wait1523;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$v37\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$v38\;
              \state\ <= pause_setI1521;
            end if;
          when pause_getII1532 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v31\ := \$arr1452_value\;
            if \$v31_lock\(0) = '1' then
              \state\ <= get_wait1530;
            else
              \$v32\ := \$v31\;
              \$v1529\ := \$arr1451_ptr_take\;
              if \$v1529\(0) = '1' then
                \state\ <= q_wait1528;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v32\));
                \state\ <= pause_getI1526;
              end if;
            end if;
          when pause_getII1536 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v30\ := \$arr1451_value\;
            \$v35\ := \$v30\(36 to 71);
            \$v1534\ := \$arr1452_ptr_take\;
            if \$v1534\(0) = '1' then
              \state\ <= q_wait1533;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1531;
            end if;
          when pause_getII1541 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v28\ := \$arr1452_value\;
            if \$v28_lock\(0) = '1' then
              \state\ <= get_wait1539;
            else
              \$v29\ := \$v28\;
              \$v1538\ := \$arr1451_ptr_take\;
              if \$v1538\(0) = '1' then
                \state\ <= q_wait1537;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v29\));
                \state\ <= pause_getI1535;
              end if;
            end if;
          when pause_getII1546 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v27\ := \$arr1452_value\;
            if \$v27_lock\(0) = '1' then
              \state\ <= get_wait1544;
            else
              \$v37\ := \$v27\;
              \$v1543\ := \$arr1452_ptr_take\;
              if \$v1543\(0) = '1' then
                \state\ <= q_wait1542;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1540;
              end if;
            end if;
          when pause_getII1554 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v24\ := \$arr1451_value\;
            \$v25\ := \$v24\(36 to 71);
            \$v1551\ := \$v25\;
            \$v1552\ := \$v1551\(0 to 3);
            \$v1550\ := \$v1551\(4 to 35);
            case \$v1552\ is
            when "0010" =>
              \$v26\ := eclat_true;
              \$v1549\ := \$v26\;
              if \$v1549\(0) = '1' then
                \$v1520\ := \$arr1452_ptr_take\;
                if \$v1520\(0) = '1' then
                  \state\ <= q_wait1519;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1517;
                end if;
              else
                \$v1548\ := \$arr1452_ptr_take\;
                if \$v1548\(0) = '1' then
                  \state\ <= q_wait1547;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1545;
                end if;
              end if;
            when others =>
              \$v26\ := eclat_false;
              \$v1549\ := \$v26\;
              if \$v1549\(0) = '1' then
                \$v1520\ := \$arr1452_ptr_take\;
                if \$v1520\(0) = '1' then
                  \state\ <= q_wait1519;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1517;
                end if;
              else
                \$v1548\ := \$arr1452_ptr_take\;
                if \$v1548\(0) = '1' then
                  \state\ <= q_wait1547;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1545;
                end if;
              end if;
            end case;
          when pause_getII1559 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v22\ := \$arr1452_value\;
            if \$v22_lock\(0) = '1' then
              \state\ <= get_wait1557;
            else
              \$v23\ := \$v22\;
              \$v1556\ := \$arr1451_ptr_take\;
              if \$v1556\(0) = '1' then
                \state\ <= q_wait1555;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v23\));
                \state\ <= pause_getI1553;
              end if;
            end if;
          when pause_getII1563 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v21\ := \$arr1451_value\;
            \$84_x\ := \$v21\(0 to 35);
            \$v1561\ := \$arr1452_ptr_take\;
            if \$v1561\(0) = '1' then
              \state\ <= q_wait1560;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1558;
            end if;
          when pause_getII1568 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v19\ := \$arr1452_value\;
            if \$v19_lock\(0) = '1' then
              \state\ <= get_wait1566;
            else
              \$v20\ := \$v19\;
              \$v1565\ := \$arr1451_ptr_take\;
              if \$v1565\(0) = '1' then
                \state\ <= q_wait1564;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v20\));
                \state\ <= pause_getI1562;
              end if;
            end if;
          when pause_getII1577 =>
            \$arr1451_ptr_take\(0) := '0';
            \$187\ := \$arr1451_value\;
            \$182\ := \$187\(36 to 71);
            \$v1574\ := \$182\;
            \$v1575\ := \$v1574\(0 to 3);
            \$v1573\ := \$v1574\(4 to 35);
            case \$v1575\ is
            when "0010" =>
              \$183_i\ := \$v1573\(0 to 31);
              \$181\ := \$183_i\;
              if \$180_lock\(0) = '1' then
                \state\ <= get_wait1571;
              else
                \$180_lock\ := eclat_true;
                \state\ <= get_pause1572;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811392\;
            end case;
          when pause_getII1582 =>
            \$arr1452_ptr_take\(0) := '0';
            \$192\ := \$arr1452_value\;
            if \$192_lock\(0) = '1' then
              \state\ <= get_wait1580;
            else
              \$191\ := \$192\;
              \$v1579\ := \$arr1451_ptr_take\;
              if \$v1579\(0) = '1' then
                \state\ <= q_wait1578;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$191\));
                \state\ <= pause_getI1576;
              end if;
            end if;
          when pause_getII1586 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1584\ := \$arr1452_ptr_take\;
            if \$v1584\(0) = '1' then
              \state\ <= q_wait1583;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1581;
            end if;
          when pause_getII1595 =>
            \$arr1451_ptr_take\(0) := '0';
            \$167\ := \$arr1451_value\;
            \$166\ := \$167\(72 to 107);
            \$v1593\ := "00000000000000000000000000000000";
            \$164\ := "0000" & \$v1593\ & \$165\ & \$166\;
            \$v1592\ := \$arr1451_ptr_take\;
            if \$v1592\(0) = '1' then
              \state\ <= q_wait1591;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$163\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$164\;
              \state\ <= pause_setI1589;
            end if;
          when pause_getII1600 =>
            \$arr1452_ptr_take\(0) := '0';
            \$172\ := \$arr1452_value\;
            if \$172_lock\(0) = '1' then
              \state\ <= get_wait1598;
            else
              \$171\ := \$172\;
              \$v1597\ := \$arr1451_ptr_take\;
              if \$v1597\(0) = '1' then
                \state\ <= q_wait1596;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$171\));
                \state\ <= pause_getI1594;
              end if;
            end if;
          when pause_getII1604 =>
            \$arr1451_ptr_take\(0) := '0';
            \$173\ := \$arr1451_value\;
            \$165\ := \$173\(36 to 71);
            \$v1602\ := \$arr1452_ptr_take\;
            if \$v1602\(0) = '1' then
              \state\ <= q_wait1601;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1599;
            end if;
          when pause_getII1609 =>
            \$arr1452_ptr_take\(0) := '0';
            \$178\ := \$arr1452_value\;
            if \$178_lock\(0) = '1' then
              \state\ <= get_wait1607;
            else
              \$177\ := \$178\;
              \$v1606\ := \$arr1451_ptr_take\;
              if \$v1606\(0) = '1' then
                \state\ <= q_wait1605;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$177\));
                \state\ <= pause_getI1603;
              end if;
            end if;
          when pause_getII1614 =>
            \$arr1452_ptr_take\(0) := '0';
            \$179\ := \$arr1452_value\;
            if \$179_lock\(0) = '1' then
              \state\ <= get_wait1612;
            else
              \$163\ := \$179\;
              \$v1611\ := \$arr1452_ptr_take\;
              if \$v1611\(0) = '1' then
                \state\ <= q_wait1610;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1608;
              end if;
            end if;
          when pause_getII1622 =>
            \$arr1451_ptr_take\(0) := '0';
            \$195\ := \$arr1451_value\;
            \$193\ := \$195\(36 to 71);
            \$v1619\ := \$193\;
            \$v1620\ := \$v1619\(0 to 3);
            \$v1618\ := \$v1619\(4 to 35);
            case \$v1620\ is
            when "0010" =>
              \$162\ := eclat_true;
              \$v1617\ := \$162\;
              if \$v1617\(0) = '1' then
                \$v1588\ := \$arr1452_ptr_take\;
                if \$v1588\(0) = '1' then
                  \state\ <= q_wait1587;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1585;
                end if;
              else
                \$v1616\ := \$arr1452_ptr_take\;
                if \$v1616\(0) = '1' then
                  \state\ <= q_wait1615;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1613;
                end if;
              end if;
            when others =>
              \$162\ := eclat_false;
              \$v1617\ := \$162\;
              if \$v1617\(0) = '1' then
                \$v1588\ := \$arr1452_ptr_take\;
                if \$v1588\(0) = '1' then
                  \state\ <= q_wait1587;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1585;
                end if;
              else
                \$v1616\ := \$arr1452_ptr_take\;
                if \$v1616\(0) = '1' then
                  \state\ <= q_wait1615;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1613;
                end if;
              end if;
            end case;
          when pause_getII1627 =>
            \$arr1452_ptr_take\(0) := '0';
            \$200\ := \$arr1452_value\;
            if \$200_lock\(0) = '1' then
              \state\ <= get_wait1625;
            else
              \$199\ := \$200\;
              \$v1624\ := \$arr1451_ptr_take\;
              if \$v1624\(0) = '1' then
                \state\ <= q_wait1623;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$199\));
                \state\ <= pause_getI1621;
              end if;
            end if;
          when pause_getII1631 =>
            \$arr1451_ptr_take\(0) := '0';
            \$201\ := \$arr1451_value\;
            \$161_x\ := \$201\(0 to 35);
            \$v1629\ := \$arr1452_ptr_take\;
            if \$v1629\(0) = '1' then
              \state\ <= q_wait1628;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1626;
            end if;
          when pause_getII1636 =>
            \$arr1452_ptr_take\(0) := '0';
            \$206\ := \$arr1452_value\;
            if \$206_lock\(0) = '1' then
              \state\ <= get_wait1634;
            else
              \$205\ := \$206\;
              \$v1633\ := \$arr1451_ptr_take\;
              if \$v1633\(0) = '1' then
                \state\ <= q_wait1632;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$205\));
                \state\ <= pause_getI1630;
              end if;
            end if;
          when pause_getII1647 =>
            \$arr1452_ptr_take\(0) := '0';
            \$219\ := \$arr1452_value\;
            if \$219_lock\(0) = '1' then
              \state\ <= get_wait1645;
            else
              \$218\ := \$219\;
              \$217\ := \$218\ & "00000000000000000000000000000001";
              \$216\ := eclat_sub(\$217\);
              if \$215_lock\(0) = '1' then
                \state\ <= get_wait1643;
              else
                \$215_lock\ := eclat_true;
                \state\ <= get_pause1644;
              end if;
            end if;
          when pause_getII1651 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1649\ := \$arr1452_ptr_take\;
            if \$v1649\(0) = '1' then
              \state\ <= q_wait1648;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1646;
            end if;
          when pause_getII1663 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$214_lock\(0) = '1' then
              \state\ <= get_wait1660;
            else
              \$214_lock\ := eclat_true;
              \state\ <= get_pause1661;
            end if;
          when pause_getII1675 =>
            \$arr1452_ptr_take\(0) := '0';
            \$220\ := \$arr1452_value\;
            if \$220_lock\(0) = '1' then
              \state\ <= get_wait1673;
            else
              \$210_i\ := \$220\;
              \$v1672\ := eclat_gt(\$210_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1672\(0) = '1' then
                \$v1671\ := eclat_eq(\$210_i\ & X"000" & X"15f90");
                if \$v1671\(0) = '1' then
                  \$v1659\ := \$arr1451_ptr_take\;
                  if \$v1659\(0) = '1' then
                    \state\ <= q_wait1658;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1654\ := "00000000000000000000000000000000";
                    \$v1655\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$209_result_after_f\ & "0001" & \$v1654\ & "0001" & \$v1655\;
                    \state\ <= pause_setI1656;
                  end if;
                else
                  \$v1670\ := \$arr1451_ptr_take\;
                  if \$v1670\(0) = '1' then
                    \state\ <= q_wait1669;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1666\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$209_result_after_f\ & "0010" & \$210_i\ & "0001" & \$v1666\;
                    \state\ <= pause_setI1667;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811393\;
              end if;
            end if;
          when pause_getII1691 =>
            \$arr1451_ptr_take\(0) := '0';
            \$250\ := \$arr1451_value\;
            \$245\ := \$250\(36 to 71);
            \$v1688\ := \$245\;
            \$v1689\ := \$v1688\(0 to 3);
            \$v1687\ := \$v1688\(4 to 35);
            case \$v1689\ is
            when "0010" =>
              \$246_i\ := \$v1687\(0 to 31);
              \$244\ := \$246_i\;
              if \$243_lock\(0) = '1' then
                \state\ <= get_wait1685;
              else
                \$243_lock\ := eclat_true;
                \state\ <= get_pause1686;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811396\;
            end case;
          when pause_getII1696 =>
            \$arr1452_ptr_take\(0) := '0';
            \$255\ := \$arr1452_value\;
            if \$255_lock\(0) = '1' then
              \state\ <= get_wait1694;
            else
              \$254\ := \$255\;
              \$v1693\ := \$arr1451_ptr_take\;
              if \$v1693\(0) = '1' then
                \state\ <= q_wait1692;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$254\));
                \state\ <= pause_getI1690;
              end if;
            end if;
          when pause_getII1700 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1698\ := \$arr1452_ptr_take\;
            if \$v1698\(0) = '1' then
              \state\ <= q_wait1697;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1695;
            end if;
          when pause_getII1709 =>
            \$arr1451_ptr_take\(0) := '0';
            \$230\ := \$arr1451_value\;
            \$229\ := \$230\(72 to 107);
            \$v1707\ := "00000000000000000000000000000000";
            \$227\ := "0000" & \$v1707\ & \$228\ & \$229\;
            \$v1706\ := \$arr1451_ptr_take\;
            if \$v1706\(0) = '1' then
              \state\ <= q_wait1705;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$226\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$227\;
              \state\ <= pause_setI1703;
            end if;
          when pause_getII1714 =>
            \$arr1452_ptr_take\(0) := '0';
            \$235\ := \$arr1452_value\;
            if \$235_lock\(0) = '1' then
              \state\ <= get_wait1712;
            else
              \$234\ := \$235\;
              \$v1711\ := \$arr1451_ptr_take\;
              if \$v1711\(0) = '1' then
                \state\ <= q_wait1710;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$234\));
                \state\ <= pause_getI1708;
              end if;
            end if;
          when pause_getII1718 =>
            \$arr1451_ptr_take\(0) := '0';
            \$236\ := \$arr1451_value\;
            \$228\ := \$236\(36 to 71);
            \$v1716\ := \$arr1452_ptr_take\;
            if \$v1716\(0) = '1' then
              \state\ <= q_wait1715;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1713;
            end if;
          when pause_getII1723 =>
            \$arr1452_ptr_take\(0) := '0';
            \$241\ := \$arr1452_value\;
            if \$241_lock\(0) = '1' then
              \state\ <= get_wait1721;
            else
              \$240\ := \$241\;
              \$v1720\ := \$arr1451_ptr_take\;
              if \$v1720\(0) = '1' then
                \state\ <= q_wait1719;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$240\));
                \state\ <= pause_getI1717;
              end if;
            end if;
          when pause_getII1728 =>
            \$arr1452_ptr_take\(0) := '0';
            \$242\ := \$arr1452_value\;
            if \$242_lock\(0) = '1' then
              \state\ <= get_wait1726;
            else
              \$226\ := \$242\;
              \$v1725\ := \$arr1452_ptr_take\;
              if \$v1725\(0) = '1' then
                \state\ <= q_wait1724;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1722;
              end if;
            end if;
          when pause_getII1736 =>
            \$arr1451_ptr_take\(0) := '0';
            \$258\ := \$arr1451_value\;
            \$256\ := \$258\(36 to 71);
            \$v1733\ := \$256\;
            \$v1734\ := \$v1733\(0 to 3);
            \$v1732\ := \$v1733\(4 to 35);
            case \$v1734\ is
            when "0010" =>
              \$225\ := eclat_true;
              \$v1731\ := \$225\;
              if \$v1731\(0) = '1' then
                \$v1702\ := \$arr1452_ptr_take\;
                if \$v1702\(0) = '1' then
                  \state\ <= q_wait1701;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1699;
                end if;
              else
                \$v1730\ := \$arr1452_ptr_take\;
                if \$v1730\(0) = '1' then
                  \state\ <= q_wait1729;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1727;
                end if;
              end if;
            when others =>
              \$225\ := eclat_false;
              \$v1731\ := \$225\;
              if \$v1731\(0) = '1' then
                \$v1702\ := \$arr1452_ptr_take\;
                if \$v1702\(0) = '1' then
                  \state\ <= q_wait1701;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1699;
                end if;
              else
                \$v1730\ := \$arr1452_ptr_take\;
                if \$v1730\(0) = '1' then
                  \state\ <= q_wait1729;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1727;
                end if;
              end if;
            end case;
          when pause_getII1741 =>
            \$arr1452_ptr_take\(0) := '0';
            \$263\ := \$arr1452_value\;
            if \$263_lock\(0) = '1' then
              \state\ <= get_wait1739;
            else
              \$262\ := \$263\;
              \$v1738\ := \$arr1451_ptr_take\;
              if \$v1738\(0) = '1' then
                \state\ <= q_wait1737;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$262\));
                \state\ <= pause_getI1735;
              end if;
            end if;
          when pause_getII1745 =>
            \$arr1451_ptr_take\(0) := '0';
            \$264\ := \$arr1451_value\;
            \$224_x\ := \$264\(0 to 35);
            \$v1743\ := \$arr1452_ptr_take\;
            if \$v1743\(0) = '1' then
              \state\ <= q_wait1742;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1740;
            end if;
          when pause_getII1750 =>
            \$arr1452_ptr_take\(0) := '0';
            \$269\ := \$arr1452_value\;
            if \$269_lock\(0) = '1' then
              \state\ <= get_wait1748;
            else
              \$268\ := \$269\;
              \$v1747\ := \$arr1451_ptr_take\;
              if \$v1747\(0) = '1' then
                \state\ <= q_wait1746;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$268\));
                \state\ <= pause_getI1744;
              end if;
            end if;
          when pause_getII1759 =>
            \$arr1451_ptr_take\(0) := '0';
            \$296\ := \$arr1451_value\;
            \$291\ := \$296\(36 to 71);
            \$v1756\ := \$291\;
            \$v1757\ := \$v1756\(0 to 3);
            \$v1755\ := \$v1756\(4 to 35);
            case \$v1757\ is
            when "0010" =>
              \$292_i\ := \$v1755\(0 to 31);
              \$290\ := \$292_i\;
              if \$289_lock\(0) = '1' then
                \state\ <= get_wait1753;
              else
                \$289_lock\ := eclat_true;
                \state\ <= get_pause1754;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811397\;
            end case;
          when pause_getII1764 =>
            \$arr1452_ptr_take\(0) := '0';
            \$301\ := \$arr1452_value\;
            if \$301_lock\(0) = '1' then
              \state\ <= get_wait1762;
            else
              \$300\ := \$301\;
              \$v1761\ := \$arr1451_ptr_take\;
              if \$v1761\(0) = '1' then
                \state\ <= q_wait1760;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$300\));
                \state\ <= pause_getI1758;
              end if;
            end if;
          when pause_getII1768 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1766\ := \$arr1452_ptr_take\;
            if \$v1766\(0) = '1' then
              \state\ <= q_wait1765;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1763;
            end if;
          when pause_getII1777 =>
            \$arr1451_ptr_take\(0) := '0';
            \$276\ := \$arr1451_value\;
            \$275\ := \$276\(72 to 107);
            \$v1775\ := "00000000000000000000000000000000";
            \$273\ := "0000" & \$v1775\ & \$274\ & \$275\;
            \$v1774\ := \$arr1451_ptr_take\;
            if \$v1774\(0) = '1' then
              \state\ <= q_wait1773;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$272\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$273\;
              \state\ <= pause_setI1771;
            end if;
          when pause_getII1782 =>
            \$arr1452_ptr_take\(0) := '0';
            \$281\ := \$arr1452_value\;
            if \$281_lock\(0) = '1' then
              \state\ <= get_wait1780;
            else
              \$280\ := \$281\;
              \$v1779\ := \$arr1451_ptr_take\;
              if \$v1779\(0) = '1' then
                \state\ <= q_wait1778;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$280\));
                \state\ <= pause_getI1776;
              end if;
            end if;
          when pause_getII1786 =>
            \$arr1451_ptr_take\(0) := '0';
            \$282\ := \$arr1451_value\;
            \$274\ := \$282\(36 to 71);
            \$v1784\ := \$arr1452_ptr_take\;
            if \$v1784\(0) = '1' then
              \state\ <= q_wait1783;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1781;
            end if;
          when pause_getII1791 =>
            \$arr1452_ptr_take\(0) := '0';
            \$287\ := \$arr1452_value\;
            if \$287_lock\(0) = '1' then
              \state\ <= get_wait1789;
            else
              \$286\ := \$287\;
              \$v1788\ := \$arr1451_ptr_take\;
              if \$v1788\(0) = '1' then
                \state\ <= q_wait1787;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$286\));
                \state\ <= pause_getI1785;
              end if;
            end if;
          when pause_getII1796 =>
            \$arr1452_ptr_take\(0) := '0';
            \$288\ := \$arr1452_value\;
            if \$288_lock\(0) = '1' then
              \state\ <= get_wait1794;
            else
              \$272\ := \$288\;
              \$v1793\ := \$arr1452_ptr_take\;
              if \$v1793\(0) = '1' then
                \state\ <= q_wait1792;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1790;
              end if;
            end if;
          when pause_getII1804 =>
            \$arr1451_ptr_take\(0) := '0';
            \$304\ := \$arr1451_value\;
            \$302\ := \$304\(36 to 71);
            \$v1801\ := \$302\;
            \$v1802\ := \$v1801\(0 to 3);
            \$v1800\ := \$v1801\(4 to 35);
            case \$v1802\ is
            when "0010" =>
              \$271\ := eclat_true;
              \$v1799\ := \$271\;
              if \$v1799\(0) = '1' then
                \$v1770\ := \$arr1452_ptr_take\;
                if \$v1770\(0) = '1' then
                  \state\ <= q_wait1769;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1767;
                end if;
              else
                \$v1798\ := \$arr1452_ptr_take\;
                if \$v1798\(0) = '1' then
                  \state\ <= q_wait1797;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1795;
                end if;
              end if;
            when others =>
              \$271\ := eclat_false;
              \$v1799\ := \$271\;
              if \$v1799\(0) = '1' then
                \$v1770\ := \$arr1452_ptr_take\;
                if \$v1770\(0) = '1' then
                  \state\ <= q_wait1769;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1767;
                end if;
              else
                \$v1798\ := \$arr1452_ptr_take\;
                if \$v1798\(0) = '1' then
                  \state\ <= q_wait1797;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1795;
                end if;
              end if;
            end case;
          when pause_getII1809 =>
            \$arr1452_ptr_take\(0) := '0';
            \$309\ := \$arr1452_value\;
            if \$309_lock\(0) = '1' then
              \state\ <= get_wait1807;
            else
              \$308\ := \$309\;
              \$v1806\ := \$arr1451_ptr_take\;
              if \$v1806\(0) = '1' then
                \state\ <= q_wait1805;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$308\));
                \state\ <= pause_getI1803;
              end if;
            end if;
          when pause_getII1813 =>
            \$arr1451_ptr_take\(0) := '0';
            \$310\ := \$arr1451_value\;
            \$270_x\ := \$310\(0 to 35);
            \$v1811\ := \$arr1452_ptr_take\;
            if \$v1811\(0) = '1' then
              \state\ <= q_wait1810;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1808;
            end if;
          when pause_getII1818 =>
            \$arr1452_ptr_take\(0) := '0';
            \$315\ := \$arr1452_value\;
            if \$315_lock\(0) = '1' then
              \state\ <= get_wait1816;
            else
              \$314\ := \$315\;
              \$v1815\ := \$arr1451_ptr_take\;
              if \$v1815\(0) = '1' then
                \state\ <= q_wait1814;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$314\));
                \state\ <= pause_getI1812;
              end if;
            end if;
          when pause_getII1829 =>
            \$arr1452_ptr_take\(0) := '0';
            \$328\ := \$arr1452_value\;
            if \$328_lock\(0) = '1' then
              \state\ <= get_wait1827;
            else
              \$327\ := \$328\;
              \$326\ := \$327\ & "00000000000000000000000000000001";
              \$325\ := eclat_sub(\$326\);
              if \$324_lock\(0) = '1' then
                \state\ <= get_wait1825;
              else
                \$324_lock\ := eclat_true;
                \state\ <= get_pause1826;
              end if;
            end if;
          when pause_getII1833 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1831\ := \$arr1452_ptr_take\;
            if \$v1831\(0) = '1' then
              \state\ <= q_wait1830;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1828;
            end if;
          when pause_getII1845 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$323_lock\(0) = '1' then
              \state\ <= get_wait1842;
            else
              \$323_lock\ := eclat_true;
              \state\ <= get_pause1843;
            end if;
          when pause_getII1857 =>
            \$arr1452_ptr_take\(0) := '0';
            \$329\ := \$arr1452_value\;
            if \$329_lock\(0) = '1' then
              \state\ <= get_wait1855;
            else
              \$319_i\ := \$329\;
              \$v1854\ := eclat_gt(\$319_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v1854\(0) = '1' then
                \$v1853\ := eclat_eq(\$319_i\ & X"000" & X"15f90");
                if \$v1853\(0) = '1' then
                  \$v1841\ := \$arr1451_ptr_take\;
                  if \$v1841\(0) = '1' then
                    \state\ <= q_wait1840;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1836\ := "00000000000000000000000000000000";
                    \$v1837\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$318_result_after_f\ & "0001" & \$v1836\ & "0001" & \$v1837\;
                    \state\ <= pause_setI1838;
                  end if;
                else
                  \$v1852\ := \$arr1451_ptr_take\;
                  if \$v1852\(0) = '1' then
                    \state\ <= q_wait1851;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v1848\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$318_result_after_f\ & "0010" & \$319_i\ & "0001" & \$v1848\;
                    \state\ <= pause_setI1849;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811398\;
              end if;
            end if;
          when pause_getII1873 =>
            \$arr1451_ptr_take\(0) := '0';
            \$359\ := \$arr1451_value\;
            \$354\ := \$359\(36 to 71);
            \$v1870\ := \$354\;
            \$v1871\ := \$v1870\(0 to 3);
            \$v1869\ := \$v1870\(4 to 35);
            case \$v1871\ is
            when "0010" =>
              \$355_i\ := \$v1869\(0 to 31);
              \$353\ := \$355_i\;
              if \$352_lock\(0) = '1' then
                \state\ <= get_wait1867;
              else
                \$352_lock\ := eclat_true;
                \state\ <= get_pause1868;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811401\;
            end case;
          when pause_getII1878 =>
            \$arr1452_ptr_take\(0) := '0';
            \$364\ := \$arr1452_value\;
            if \$364_lock\(0) = '1' then
              \state\ <= get_wait1876;
            else
              \$363\ := \$364\;
              \$v1875\ := \$arr1451_ptr_take\;
              if \$v1875\(0) = '1' then
                \state\ <= q_wait1874;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$363\));
                \state\ <= pause_getI1872;
              end if;
            end if;
          when pause_getII1882 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1880\ := \$arr1452_ptr_take\;
            if \$v1880\(0) = '1' then
              \state\ <= q_wait1879;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1877;
            end if;
          when pause_getII1891 =>
            \$arr1451_ptr_take\(0) := '0';
            \$339\ := \$arr1451_value\;
            \$338\ := \$339\(72 to 107);
            \$v1889\ := "00000000000000000000000000000000";
            \$336\ := "0000" & \$v1889\ & \$337\ & \$338\;
            \$v1888\ := \$arr1451_ptr_take\;
            if \$v1888\(0) = '1' then
              \state\ <= q_wait1887;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$335\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$336\;
              \state\ <= pause_setI1885;
            end if;
          when pause_getII1896 =>
            \$arr1452_ptr_take\(0) := '0';
            \$344\ := \$arr1452_value\;
            if \$344_lock\(0) = '1' then
              \state\ <= get_wait1894;
            else
              \$343\ := \$344\;
              \$v1893\ := \$arr1451_ptr_take\;
              if \$v1893\(0) = '1' then
                \state\ <= q_wait1892;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$343\));
                \state\ <= pause_getI1890;
              end if;
            end if;
          when pause_getII1900 =>
            \$arr1451_ptr_take\(0) := '0';
            \$345\ := \$arr1451_value\;
            \$337\ := \$345\(36 to 71);
            \$v1898\ := \$arr1452_ptr_take\;
            if \$v1898\(0) = '1' then
              \state\ <= q_wait1897;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1895;
            end if;
          when pause_getII1905 =>
            \$arr1452_ptr_take\(0) := '0';
            \$350\ := \$arr1452_value\;
            if \$350_lock\(0) = '1' then
              \state\ <= get_wait1903;
            else
              \$349\ := \$350\;
              \$v1902\ := \$arr1451_ptr_take\;
              if \$v1902\(0) = '1' then
                \state\ <= q_wait1901;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$349\));
                \state\ <= pause_getI1899;
              end if;
            end if;
          when pause_getII1910 =>
            \$arr1452_ptr_take\(0) := '0';
            \$351\ := \$arr1452_value\;
            if \$351_lock\(0) = '1' then
              \state\ <= get_wait1908;
            else
              \$335\ := \$351\;
              \$v1907\ := \$arr1452_ptr_take\;
              if \$v1907\(0) = '1' then
                \state\ <= q_wait1906;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1904;
              end if;
            end if;
          when pause_getII1918 =>
            \$arr1451_ptr_take\(0) := '0';
            \$367\ := \$arr1451_value\;
            \$365\ := \$367\(36 to 71);
            \$v1915\ := \$365\;
            \$v1916\ := \$v1915\(0 to 3);
            \$v1914\ := \$v1915\(4 to 35);
            case \$v1916\ is
            when "0010" =>
              \$334\ := eclat_true;
              \$v1913\ := \$334\;
              if \$v1913\(0) = '1' then
                \$v1884\ := \$arr1452_ptr_take\;
                if \$v1884\(0) = '1' then
                  \state\ <= q_wait1883;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1881;
                end if;
              else
                \$v1912\ := \$arr1452_ptr_take\;
                if \$v1912\(0) = '1' then
                  \state\ <= q_wait1911;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1909;
                end if;
              end if;
            when others =>
              \$334\ := eclat_false;
              \$v1913\ := \$334\;
              if \$v1913\(0) = '1' then
                \$v1884\ := \$arr1452_ptr_take\;
                if \$v1884\(0) = '1' then
                  \state\ <= q_wait1883;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1881;
                end if;
              else
                \$v1912\ := \$arr1452_ptr_take\;
                if \$v1912\(0) = '1' then
                  \state\ <= q_wait1911;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1909;
                end if;
              end if;
            end case;
          when pause_getII1923 =>
            \$arr1452_ptr_take\(0) := '0';
            \$372\ := \$arr1452_value\;
            if \$372_lock\(0) = '1' then
              \state\ <= get_wait1921;
            else
              \$371\ := \$372\;
              \$v1920\ := \$arr1451_ptr_take\;
              if \$v1920\(0) = '1' then
                \state\ <= q_wait1919;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$371\));
                \state\ <= pause_getI1917;
              end if;
            end if;
          when pause_getII1927 =>
            \$arr1451_ptr_take\(0) := '0';
            \$373\ := \$arr1451_value\;
            \$333_x\ := \$373\(0 to 35);
            \$v1925\ := \$arr1452_ptr_take\;
            if \$v1925\(0) = '1' then
              \state\ <= q_wait1924;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1922;
            end if;
          when pause_getII1932 =>
            \$arr1452_ptr_take\(0) := '0';
            \$378\ := \$arr1452_value\;
            if \$378_lock\(0) = '1' then
              \state\ <= get_wait1930;
            else
              \$377\ := \$378\;
              \$v1929\ := \$arr1451_ptr_take\;
              if \$v1929\(0) = '1' then
                \state\ <= q_wait1928;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$377\));
                \state\ <= pause_getI1926;
              end if;
            end if;
          when pause_getII1941 =>
            \$arr1451_ptr_take\(0) := '0';
            \$405\ := \$arr1451_value\;
            \$400\ := \$405\(36 to 71);
            \$v1938\ := \$400\;
            \$v1939\ := \$v1938\(0 to 3);
            \$v1937\ := \$v1938\(4 to 35);
            case \$v1939\ is
            when "0010" =>
              \$401_i\ := \$v1937\(0 to 31);
              \$399\ := \$401_i\;
              if \$398_lock\(0) = '1' then
                \state\ <= get_wait1935;
              else
                \$398_lock\ := eclat_true;
                \state\ <= get_pause1936;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811402\;
            end case;
          when pause_getII1946 =>
            \$arr1452_ptr_take\(0) := '0';
            \$410\ := \$arr1452_value\;
            if \$410_lock\(0) = '1' then
              \state\ <= get_wait1944;
            else
              \$409\ := \$410\;
              \$v1943\ := \$arr1451_ptr_take\;
              if \$v1943\(0) = '1' then
                \state\ <= q_wait1942;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$409\));
                \state\ <= pause_getI1940;
              end if;
            end if;
          when pause_getII1950 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v1948\ := \$arr1452_ptr_take\;
            if \$v1948\(0) = '1' then
              \state\ <= q_wait1947;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1945;
            end if;
          when pause_getII1959 =>
            \$arr1451_ptr_take\(0) := '0';
            \$385\ := \$arr1451_value\;
            \$384\ := \$385\(72 to 107);
            \$v1957\ := "00000000000000000000000000000000";
            \$382\ := "0000" & \$v1957\ & \$383\ & \$384\;
            \$v1956\ := \$arr1451_ptr_take\;
            if \$v1956\(0) = '1' then
              \state\ <= q_wait1955;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$381\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$382\;
              \state\ <= pause_setI1953;
            end if;
          when pause_getII1964 =>
            \$arr1452_ptr_take\(0) := '0';
            \$390\ := \$arr1452_value\;
            if \$390_lock\(0) = '1' then
              \state\ <= get_wait1962;
            else
              \$389\ := \$390\;
              \$v1961\ := \$arr1451_ptr_take\;
              if \$v1961\(0) = '1' then
                \state\ <= q_wait1960;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$389\));
                \state\ <= pause_getI1958;
              end if;
            end if;
          when pause_getII1968 =>
            \$arr1451_ptr_take\(0) := '0';
            \$391\ := \$arr1451_value\;
            \$383\ := \$391\(36 to 71);
            \$v1966\ := \$arr1452_ptr_take\;
            if \$v1966\(0) = '1' then
              \state\ <= q_wait1965;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1963;
            end if;
          when pause_getII1973 =>
            \$arr1452_ptr_take\(0) := '0';
            \$396\ := \$arr1452_value\;
            if \$396_lock\(0) = '1' then
              \state\ <= get_wait1971;
            else
              \$395\ := \$396\;
              \$v1970\ := \$arr1451_ptr_take\;
              if \$v1970\(0) = '1' then
                \state\ <= q_wait1969;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$395\));
                \state\ <= pause_getI1967;
              end if;
            end if;
          when pause_getII1978 =>
            \$arr1452_ptr_take\(0) := '0';
            \$397\ := \$arr1452_value\;
            if \$397_lock\(0) = '1' then
              \state\ <= get_wait1976;
            else
              \$381\ := \$397\;
              \$v1975\ := \$arr1452_ptr_take\;
              if \$v1975\(0) = '1' then
                \state\ <= q_wait1974;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI1972;
              end if;
            end if;
          when pause_getII1986 =>
            \$arr1451_ptr_take\(0) := '0';
            \$413\ := \$arr1451_value\;
            \$411\ := \$413\(36 to 71);
            \$v1983\ := \$411\;
            \$v1984\ := \$v1983\(0 to 3);
            \$v1982\ := \$v1983\(4 to 35);
            case \$v1984\ is
            when "0010" =>
              \$380\ := eclat_true;
              \$v1981\ := \$380\;
              if \$v1981\(0) = '1' then
                \$v1952\ := \$arr1452_ptr_take\;
                if \$v1952\(0) = '1' then
                  \state\ <= q_wait1951;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1949;
                end if;
              else
                \$v1980\ := \$arr1452_ptr_take\;
                if \$v1980\(0) = '1' then
                  \state\ <= q_wait1979;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1977;
                end if;
              end if;
            when others =>
              \$380\ := eclat_false;
              \$v1981\ := \$380\;
              if \$v1981\(0) = '1' then
                \$v1952\ := \$arr1452_ptr_take\;
                if \$v1952\(0) = '1' then
                  \state\ <= q_wait1951;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1949;
                end if;
              else
                \$v1980\ := \$arr1452_ptr_take\;
                if \$v1980\(0) = '1' then
                  \state\ <= q_wait1979;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1977;
                end if;
              end if;
            end case;
          when pause_getII1991 =>
            \$arr1452_ptr_take\(0) := '0';
            \$418\ := \$arr1452_value\;
            if \$418_lock\(0) = '1' then
              \state\ <= get_wait1989;
            else
              \$417\ := \$418\;
              \$v1988\ := \$arr1451_ptr_take\;
              if \$v1988\(0) = '1' then
                \state\ <= q_wait1987;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$417\));
                \state\ <= pause_getI1985;
              end if;
            end if;
          when pause_getII1995 =>
            \$arr1451_ptr_take\(0) := '0';
            \$419\ := \$arr1451_value\;
            \$379_x\ := \$419\(0 to 35);
            \$v1993\ := \$arr1452_ptr_take\;
            if \$v1993\(0) = '1' then
              \state\ <= q_wait1992;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1990;
            end if;
          when pause_getII2000 =>
            \$arr1452_ptr_take\(0) := '0';
            \$424\ := \$arr1452_value\;
            if \$424_lock\(0) = '1' then
              \state\ <= get_wait1998;
            else
              \$423\ := \$424\;
              \$v1997\ := \$arr1451_ptr_take\;
              if \$v1997\(0) = '1' then
                \state\ <= q_wait1996;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$423\));
                \state\ <= pause_getI1994;
              end if;
            end if;
          when pause_getII2011 =>
            \$arr1452_ptr_take\(0) := '0';
            \$437\ := \$arr1452_value\;
            if \$437_lock\(0) = '1' then
              \state\ <= get_wait2009;
            else
              \$436\ := \$437\;
              \$435\ := \$436\ & "00000000000000000000000000000001";
              \$434\ := eclat_sub(\$435\);
              if \$433_lock\(0) = '1' then
                \state\ <= get_wait2007;
              else
                \$433_lock\ := eclat_true;
                \state\ <= get_pause2008;
              end if;
            end if;
          when pause_getII2015 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2013\ := \$arr1452_ptr_take\;
            if \$v2013\(0) = '1' then
              \state\ <= q_wait2012;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2010;
            end if;
          when pause_getII2027 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$432_lock\(0) = '1' then
              \state\ <= get_wait2024;
            else
              \$432_lock\ := eclat_true;
              \state\ <= get_pause2025;
            end if;
          when pause_getII2039 =>
            \$arr1452_ptr_take\(0) := '0';
            \$438\ := \$arr1452_value\;
            if \$438_lock\(0) = '1' then
              \state\ <= get_wait2037;
            else
              \$428_i\ := \$438\;
              \$v2036\ := eclat_gt(\$428_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2036\(0) = '1' then
                \$v2035\ := eclat_eq(\$428_i\ & X"000" & X"15f90");
                if \$v2035\(0) = '1' then
                  \$v2023\ := \$arr1451_ptr_take\;
                  if \$v2023\(0) = '1' then
                    \state\ <= q_wait2022;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2018\ := "00000000000000000000000000000000";
                    \$v2019\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$427_result_after_f\ & "0001" & \$v2018\ & "0001" & \$v2019\;
                    \state\ <= pause_setI2020;
                  end if;
                else
                  \$v2034\ := \$arr1451_ptr_take\;
                  if \$v2034\(0) = '1' then
                    \state\ <= q_wait2033;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2030\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$427_result_after_f\ & "0010" & \$428_i\ & "0001" & \$v2030\;
                    \state\ <= pause_setI2031;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811403\;
              end if;
            end if;
          when pause_getII2055 =>
            \$arr1451_ptr_take\(0) := '0';
            \$468\ := \$arr1451_value\;
            \$463\ := \$468\(36 to 71);
            \$v2052\ := \$463\;
            \$v2053\ := \$v2052\(0 to 3);
            \$v2051\ := \$v2052\(4 to 35);
            case \$v2053\ is
            when "0010" =>
              \$464_i\ := \$v2051\(0 to 31);
              \$462\ := \$464_i\;
              if \$461_lock\(0) = '1' then
                \state\ <= get_wait2049;
              else
                \$461_lock\ := eclat_true;
                \state\ <= get_pause2050;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811406\;
            end case;
          when pause_getII2060 =>
            \$arr1452_ptr_take\(0) := '0';
            \$473\ := \$arr1452_value\;
            if \$473_lock\(0) = '1' then
              \state\ <= get_wait2058;
            else
              \$472\ := \$473\;
              \$v2057\ := \$arr1451_ptr_take\;
              if \$v2057\(0) = '1' then
                \state\ <= q_wait2056;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$472\));
                \state\ <= pause_getI2054;
              end if;
            end if;
          when pause_getII2064 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2062\ := \$arr1452_ptr_take\;
            if \$v2062\(0) = '1' then
              \state\ <= q_wait2061;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2059;
            end if;
          when pause_getII2073 =>
            \$arr1451_ptr_take\(0) := '0';
            \$448\ := \$arr1451_value\;
            \$447\ := \$448\(72 to 107);
            \$v2071\ := "00000000000000000000000000000000";
            \$445\ := "0000" & \$v2071\ & \$446\ & \$447\;
            \$v2070\ := \$arr1451_ptr_take\;
            if \$v2070\(0) = '1' then
              \state\ <= q_wait2069;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$444\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$445\;
              \state\ <= pause_setI2067;
            end if;
          when pause_getII2078 =>
            \$arr1452_ptr_take\(0) := '0';
            \$453\ := \$arr1452_value\;
            if \$453_lock\(0) = '1' then
              \state\ <= get_wait2076;
            else
              \$452\ := \$453\;
              \$v2075\ := \$arr1451_ptr_take\;
              if \$v2075\(0) = '1' then
                \state\ <= q_wait2074;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$452\));
                \state\ <= pause_getI2072;
              end if;
            end if;
          when pause_getII2082 =>
            \$arr1451_ptr_take\(0) := '0';
            \$454\ := \$arr1451_value\;
            \$446\ := \$454\(36 to 71);
            \$v2080\ := \$arr1452_ptr_take\;
            if \$v2080\(0) = '1' then
              \state\ <= q_wait2079;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2077;
            end if;
          when pause_getII2087 =>
            \$arr1452_ptr_take\(0) := '0';
            \$459\ := \$arr1452_value\;
            if \$459_lock\(0) = '1' then
              \state\ <= get_wait2085;
            else
              \$458\ := \$459\;
              \$v2084\ := \$arr1451_ptr_take\;
              if \$v2084\(0) = '1' then
                \state\ <= q_wait2083;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$458\));
                \state\ <= pause_getI2081;
              end if;
            end if;
          when pause_getII2092 =>
            \$arr1452_ptr_take\(0) := '0';
            \$460\ := \$arr1452_value\;
            if \$460_lock\(0) = '1' then
              \state\ <= get_wait2090;
            else
              \$444\ := \$460\;
              \$v2089\ := \$arr1452_ptr_take\;
              if \$v2089\(0) = '1' then
                \state\ <= q_wait2088;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2086;
              end if;
            end if;
          when pause_getII2100 =>
            \$arr1451_ptr_take\(0) := '0';
            \$476\ := \$arr1451_value\;
            \$474\ := \$476\(36 to 71);
            \$v2097\ := \$474\;
            \$v2098\ := \$v2097\(0 to 3);
            \$v2096\ := \$v2097\(4 to 35);
            case \$v2098\ is
            when "0010" =>
              \$443\ := eclat_true;
              \$v2095\ := \$443\;
              if \$v2095\(0) = '1' then
                \$v2066\ := \$arr1452_ptr_take\;
                if \$v2066\(0) = '1' then
                  \state\ <= q_wait2065;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2063;
                end if;
              else
                \$v2094\ := \$arr1452_ptr_take\;
                if \$v2094\(0) = '1' then
                  \state\ <= q_wait2093;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2091;
                end if;
              end if;
            when others =>
              \$443\ := eclat_false;
              \$v2095\ := \$443\;
              if \$v2095\(0) = '1' then
                \$v2066\ := \$arr1452_ptr_take\;
                if \$v2066\(0) = '1' then
                  \state\ <= q_wait2065;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2063;
                end if;
              else
                \$v2094\ := \$arr1452_ptr_take\;
                if \$v2094\(0) = '1' then
                  \state\ <= q_wait2093;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2091;
                end if;
              end if;
            end case;
          when pause_getII2105 =>
            \$arr1452_ptr_take\(0) := '0';
            \$481\ := \$arr1452_value\;
            if \$481_lock\(0) = '1' then
              \state\ <= get_wait2103;
            else
              \$480\ := \$481\;
              \$v2102\ := \$arr1451_ptr_take\;
              if \$v2102\(0) = '1' then
                \state\ <= q_wait2101;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$480\));
                \state\ <= pause_getI2099;
              end if;
            end if;
          when pause_getII2109 =>
            \$arr1451_ptr_take\(0) := '0';
            \$482\ := \$arr1451_value\;
            \$442_x\ := \$482\(0 to 35);
            \$v2107\ := \$arr1452_ptr_take\;
            if \$v2107\(0) = '1' then
              \state\ <= q_wait2106;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2104;
            end if;
          when pause_getII2114 =>
            \$arr1452_ptr_take\(0) := '0';
            \$487\ := \$arr1452_value\;
            if \$487_lock\(0) = '1' then
              \state\ <= get_wait2112;
            else
              \$486\ := \$487\;
              \$v2111\ := \$arr1451_ptr_take\;
              if \$v2111\(0) = '1' then
                \state\ <= q_wait2110;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$486\));
                \state\ <= pause_getI2108;
              end if;
            end if;
          when pause_getII2123 =>
            \$arr1451_ptr_take\(0) := '0';
            \$514\ := \$arr1451_value\;
            \$509\ := \$514\(36 to 71);
            \$v2120\ := \$509\;
            \$v2121\ := \$v2120\(0 to 3);
            \$v2119\ := \$v2120\(4 to 35);
            case \$v2121\ is
            when "0010" =>
              \$510_i\ := \$v2119\(0 to 31);
              \$508\ := \$510_i\;
              if \$507_lock\(0) = '1' then
                \state\ <= get_wait2117;
              else
                \$507_lock\ := eclat_true;
                \state\ <= get_pause2118;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811407\;
            end case;
          when pause_getII2128 =>
            \$arr1452_ptr_take\(0) := '0';
            \$519\ := \$arr1452_value\;
            if \$519_lock\(0) = '1' then
              \state\ <= get_wait2126;
            else
              \$518\ := \$519\;
              \$v2125\ := \$arr1451_ptr_take\;
              if \$v2125\(0) = '1' then
                \state\ <= q_wait2124;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$518\));
                \state\ <= pause_getI2122;
              end if;
            end if;
          when pause_getII2132 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2130\ := \$arr1452_ptr_take\;
            if \$v2130\(0) = '1' then
              \state\ <= q_wait2129;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2127;
            end if;
          when pause_getII2141 =>
            \$arr1451_ptr_take\(0) := '0';
            \$494\ := \$arr1451_value\;
            \$493\ := \$494\(72 to 107);
            \$v2139\ := "00000000000000000000000000000000";
            \$491\ := "0000" & \$v2139\ & \$492\ & \$493\;
            \$v2138\ := \$arr1451_ptr_take\;
            if \$v2138\(0) = '1' then
              \state\ <= q_wait2137;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$490\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$491\;
              \state\ <= pause_setI2135;
            end if;
          when pause_getII2146 =>
            \$arr1452_ptr_take\(0) := '0';
            \$499\ := \$arr1452_value\;
            if \$499_lock\(0) = '1' then
              \state\ <= get_wait2144;
            else
              \$498\ := \$499\;
              \$v2143\ := \$arr1451_ptr_take\;
              if \$v2143\(0) = '1' then
                \state\ <= q_wait2142;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$498\));
                \state\ <= pause_getI2140;
              end if;
            end if;
          when pause_getII2150 =>
            \$arr1451_ptr_take\(0) := '0';
            \$500\ := \$arr1451_value\;
            \$492\ := \$500\(36 to 71);
            \$v2148\ := \$arr1452_ptr_take\;
            if \$v2148\(0) = '1' then
              \state\ <= q_wait2147;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2145;
            end if;
          when pause_getII2155 =>
            \$arr1452_ptr_take\(0) := '0';
            \$505\ := \$arr1452_value\;
            if \$505_lock\(0) = '1' then
              \state\ <= get_wait2153;
            else
              \$504\ := \$505\;
              \$v2152\ := \$arr1451_ptr_take\;
              if \$v2152\(0) = '1' then
                \state\ <= q_wait2151;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$504\));
                \state\ <= pause_getI2149;
              end if;
            end if;
          when pause_getII2160 =>
            \$arr1452_ptr_take\(0) := '0';
            \$506\ := \$arr1452_value\;
            if \$506_lock\(0) = '1' then
              \state\ <= get_wait2158;
            else
              \$490\ := \$506\;
              \$v2157\ := \$arr1452_ptr_take\;
              if \$v2157\(0) = '1' then
                \state\ <= q_wait2156;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2154;
              end if;
            end if;
          when pause_getII2168 =>
            \$arr1451_ptr_take\(0) := '0';
            \$522\ := \$arr1451_value\;
            \$520\ := \$522\(36 to 71);
            \$v2165\ := \$520\;
            \$v2166\ := \$v2165\(0 to 3);
            \$v2164\ := \$v2165\(4 to 35);
            case \$v2166\ is
            when "0010" =>
              \$489\ := eclat_true;
              \$v2163\ := \$489\;
              if \$v2163\(0) = '1' then
                \$v2134\ := \$arr1452_ptr_take\;
                if \$v2134\(0) = '1' then
                  \state\ <= q_wait2133;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2131;
                end if;
              else
                \$v2162\ := \$arr1452_ptr_take\;
                if \$v2162\(0) = '1' then
                  \state\ <= q_wait2161;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2159;
                end if;
              end if;
            when others =>
              \$489\ := eclat_false;
              \$v2163\ := \$489\;
              if \$v2163\(0) = '1' then
                \$v2134\ := \$arr1452_ptr_take\;
                if \$v2134\(0) = '1' then
                  \state\ <= q_wait2133;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2131;
                end if;
              else
                \$v2162\ := \$arr1452_ptr_take\;
                if \$v2162\(0) = '1' then
                  \state\ <= q_wait2161;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2159;
                end if;
              end if;
            end case;
          when pause_getII2173 =>
            \$arr1452_ptr_take\(0) := '0';
            \$527\ := \$arr1452_value\;
            if \$527_lock\(0) = '1' then
              \state\ <= get_wait2171;
            else
              \$526\ := \$527\;
              \$v2170\ := \$arr1451_ptr_take\;
              if \$v2170\(0) = '1' then
                \state\ <= q_wait2169;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$526\));
                \state\ <= pause_getI2167;
              end if;
            end if;
          when pause_getII2177 =>
            \$arr1451_ptr_take\(0) := '0';
            \$528\ := \$arr1451_value\;
            \$488_x\ := \$528\(0 to 35);
            \$v2175\ := \$arr1452_ptr_take\;
            if \$v2175\(0) = '1' then
              \state\ <= q_wait2174;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2172;
            end if;
          when pause_getII2182 =>
            \$arr1452_ptr_take\(0) := '0';
            \$533\ := \$arr1452_value\;
            if \$533_lock\(0) = '1' then
              \state\ <= get_wait2180;
            else
              \$532\ := \$533\;
              \$v2179\ := \$arr1451_ptr_take\;
              if \$v2179\(0) = '1' then
                \state\ <= q_wait2178;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$532\));
                \state\ <= pause_getI2176;
              end if;
            end if;
          when pause_getII2192 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$v58_lock\(0) = '1' then
              \state\ <= get_wait2189;
            else
              \$v58_lock\ := eclat_true;
              \state\ <= get_pause2190;
            end if;
          when pause_getII2208 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$v55_lock\(0) = '1' then
              \state\ <= get_wait2205;
            else
              \$v55_lock\ := eclat_true;
              \state\ <= get_pause2206;
            end if;
          when pause_getII2231 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v45\ := \$arr1452_value\;
            if \$v45_lock\(0) = '1' then
              \state\ <= get_wait2229;
            else
              \$82_i\ := \$v45\;
              \$v2228\ := eclat_gt(\$82_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2228\(0) = '1' then
                \$v2227\ := eclat_eq(\$82_i\ & X"000" & X"15f90");
                if \$v2227\(0) = '1' then
                  \$v2204\ := \$arr1451_ptr_take\;
                  if \$v2204\(0) = '1' then
                    \state\ <= q_wait2203;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2198\ := "00000000000000000000000000000000";
                    \$v2199\ := "00000000000000000000000000000000";
                    \$v2200\ := "00000000000000000000000000000101";
                    \$v2195\ := "00000000000000000000000000000000";
                    \$v2196\ := "00000000000000000000000000000000";
                    \$v2197\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(result & "0001" & \$v2198\ & "0001" & \$v2199\ & "0001" & \$v2200\ & "0001" & \$v2195\ & "0001" & \$v2196\ & "0001" & \$v2197\);
                    \state\ <= pause_setI2201;
                  end if;
                else
                  \$v2226\ := \$arr1451_ptr_take\;
                  if \$v2226\(0) = '1' then
                    \state\ <= q_wait2225;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2220\ := "00000000000000000000000000000000";
                    \$v2221\ := "00000000000000000000000000000000";
                    \$v2222\ := "00000000000000000000000000000101";
                    \$v2217\ := "00000000000000000000000000000000";
                    \$v2218\ := "00000000000000000000000000000000";
                    \$v2219\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(result & "0001" & \$v2220\ & "0001" & \$v2221\ & "0001" & \$v2222\ & "0001" & \$v2217\ & "0001" & \$v2218\ & "0001" & \$v2219\);
                    \state\ <= pause_setI2223;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811408\;
              end if;
            end if;
          when pause_getII2246 =>
            \$arr1451_ptr_take\(0) := '0';
            \$566\ := \$arr1451_value\;
            \$561\ := \$566\(36 to 71);
            \$v2243\ := \$561\;
            \$v2244\ := \$v2243\(0 to 3);
            \$v2242\ := \$v2243\(4 to 35);
            case \$v2244\ is
            when "0010" =>
              \$562_i\ := \$v2242\(0 to 31);
              \$560\ := \$562_i\;
              if \$559_lock\(0) = '1' then
                \state\ <= get_wait2240;
              else
                \$559_lock\ := eclat_true;
                \state\ <= get_pause2241;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811411\;
            end case;
          when pause_getII2251 =>
            \$arr1452_ptr_take\(0) := '0';
            \$571\ := \$arr1452_value\;
            if \$571_lock\(0) = '1' then
              \state\ <= get_wait2249;
            else
              \$570\ := \$571\;
              \$v2248\ := \$arr1451_ptr_take\;
              if \$v2248\(0) = '1' then
                \state\ <= q_wait2247;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$570\));
                \state\ <= pause_getI2245;
              end if;
            end if;
          when pause_getII2255 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2253\ := \$arr1452_ptr_take\;
            if \$v2253\(0) = '1' then
              \state\ <= q_wait2252;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2250;
            end if;
          when pause_getII2264 =>
            \$arr1451_ptr_take\(0) := '0';
            \$546\ := \$arr1451_value\;
            \$545\ := \$546\(72 to 107);
            \$v2262\ := "00000000000000000000000000000000";
            \$543\ := "0000" & \$v2262\ & \$544\ & \$545\;
            \$v2261\ := \$arr1451_ptr_take\;
            if \$v2261\(0) = '1' then
              \state\ <= q_wait2260;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$542\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$543\;
              \state\ <= pause_setI2258;
            end if;
          when pause_getII2269 =>
            \$arr1452_ptr_take\(0) := '0';
            \$551\ := \$arr1452_value\;
            if \$551_lock\(0) = '1' then
              \state\ <= get_wait2267;
            else
              \$550\ := \$551\;
              \$v2266\ := \$arr1451_ptr_take\;
              if \$v2266\(0) = '1' then
                \state\ <= q_wait2265;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$550\));
                \state\ <= pause_getI2263;
              end if;
            end if;
          when pause_getII2273 =>
            \$arr1451_ptr_take\(0) := '0';
            \$552\ := \$arr1451_value\;
            \$544\ := \$552\(36 to 71);
            \$v2271\ := \$arr1452_ptr_take\;
            if \$v2271\(0) = '1' then
              \state\ <= q_wait2270;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2268;
            end if;
          when pause_getII2278 =>
            \$arr1452_ptr_take\(0) := '0';
            \$557\ := \$arr1452_value\;
            if \$557_lock\(0) = '1' then
              \state\ <= get_wait2276;
            else
              \$556\ := \$557\;
              \$v2275\ := \$arr1451_ptr_take\;
              if \$v2275\(0) = '1' then
                \state\ <= q_wait2274;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$556\));
                \state\ <= pause_getI2272;
              end if;
            end if;
          when pause_getII2283 =>
            \$arr1452_ptr_take\(0) := '0';
            \$558\ := \$arr1452_value\;
            if \$558_lock\(0) = '1' then
              \state\ <= get_wait2281;
            else
              \$542\ := \$558\;
              \$v2280\ := \$arr1452_ptr_take\;
              if \$v2280\(0) = '1' then
                \state\ <= q_wait2279;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2277;
              end if;
            end if;
          when pause_getII2291 =>
            \$arr1451_ptr_take\(0) := '0';
            \$574\ := \$arr1451_value\;
            \$572\ := \$574\(36 to 71);
            \$v2288\ := \$572\;
            \$v2289\ := \$v2288\(0 to 3);
            \$v2287\ := \$v2288\(4 to 35);
            case \$v2289\ is
            when "0010" =>
              \$541\ := eclat_true;
              \$v2286\ := \$541\;
              if \$v2286\(0) = '1' then
                \$v2257\ := \$arr1452_ptr_take\;
                if \$v2257\(0) = '1' then
                  \state\ <= q_wait2256;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2254;
                end if;
              else
                \$v2285\ := \$arr1452_ptr_take\;
                if \$v2285\(0) = '1' then
                  \state\ <= q_wait2284;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2282;
                end if;
              end if;
            when others =>
              \$541\ := eclat_false;
              \$v2286\ := \$541\;
              if \$v2286\(0) = '1' then
                \$v2257\ := \$arr1452_ptr_take\;
                if \$v2257\(0) = '1' then
                  \state\ <= q_wait2256;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2254;
                end if;
              else
                \$v2285\ := \$arr1452_ptr_take\;
                if \$v2285\(0) = '1' then
                  \state\ <= q_wait2284;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2282;
                end if;
              end if;
            end case;
          when pause_getII2296 =>
            \$arr1452_ptr_take\(0) := '0';
            \$579\ := \$arr1452_value\;
            if \$579_lock\(0) = '1' then
              \state\ <= get_wait2294;
            else
              \$578\ := \$579\;
              \$v2293\ := \$arr1451_ptr_take\;
              if \$v2293\(0) = '1' then
                \state\ <= q_wait2292;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$578\));
                \state\ <= pause_getI2290;
              end if;
            end if;
          when pause_getII2300 =>
            \$arr1451_ptr_take\(0) := '0';
            \$580\ := \$arr1451_value\;
            \$540_x\ := \$580\(0 to 35);
            \$v2298\ := \$arr1452_ptr_take\;
            if \$v2298\(0) = '1' then
              \state\ <= q_wait2297;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2295;
            end if;
          when pause_getII2305 =>
            \$arr1452_ptr_take\(0) := '0';
            \$585\ := \$arr1452_value\;
            if \$585_lock\(0) = '1' then
              \state\ <= get_wait2303;
            else
              \$584\ := \$585\;
              \$v2302\ := \$arr1451_ptr_take\;
              if \$v2302\(0) = '1' then
                \state\ <= q_wait2301;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$584\));
                \state\ <= pause_getI2299;
              end if;
            end if;
          when pause_getII2314 =>
            \$arr1451_ptr_take\(0) := '0';
            \$612\ := \$arr1451_value\;
            \$607\ := \$612\(36 to 71);
            \$v2311\ := \$607\;
            \$v2312\ := \$v2311\(0 to 3);
            \$v2310\ := \$v2311\(4 to 35);
            case \$v2312\ is
            when "0010" =>
              \$608_i\ := \$v2310\(0 to 31);
              \$606\ := \$608_i\;
              if \$605_lock\(0) = '1' then
                \state\ <= get_wait2308;
              else
                \$605_lock\ := eclat_true;
                \state\ <= get_pause2309;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811412\;
            end case;
          when pause_getII2319 =>
            \$arr1452_ptr_take\(0) := '0';
            \$617\ := \$arr1452_value\;
            if \$617_lock\(0) = '1' then
              \state\ <= get_wait2317;
            else
              \$616\ := \$617\;
              \$v2316\ := \$arr1451_ptr_take\;
              if \$v2316\(0) = '1' then
                \state\ <= q_wait2315;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$616\));
                \state\ <= pause_getI2313;
              end if;
            end if;
          when pause_getII2323 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2321\ := \$arr1452_ptr_take\;
            if \$v2321\(0) = '1' then
              \state\ <= q_wait2320;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2318;
            end if;
          when pause_getII2332 =>
            \$arr1451_ptr_take\(0) := '0';
            \$592\ := \$arr1451_value\;
            \$591\ := \$592\(72 to 107);
            \$v2330\ := "00000000000000000000000000000000";
            \$589\ := "0000" & \$v2330\ & \$590\ & \$591\;
            \$v2329\ := \$arr1451_ptr_take\;
            if \$v2329\(0) = '1' then
              \state\ <= q_wait2328;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$588\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$589\;
              \state\ <= pause_setI2326;
            end if;
          when pause_getII2337 =>
            \$arr1452_ptr_take\(0) := '0';
            \$597\ := \$arr1452_value\;
            if \$597_lock\(0) = '1' then
              \state\ <= get_wait2335;
            else
              \$596\ := \$597\;
              \$v2334\ := \$arr1451_ptr_take\;
              if \$v2334\(0) = '1' then
                \state\ <= q_wait2333;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$596\));
                \state\ <= pause_getI2331;
              end if;
            end if;
          when pause_getII2341 =>
            \$arr1451_ptr_take\(0) := '0';
            \$598\ := \$arr1451_value\;
            \$590\ := \$598\(36 to 71);
            \$v2339\ := \$arr1452_ptr_take\;
            if \$v2339\(0) = '1' then
              \state\ <= q_wait2338;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2336;
            end if;
          when pause_getII2346 =>
            \$arr1452_ptr_take\(0) := '0';
            \$603\ := \$arr1452_value\;
            if \$603_lock\(0) = '1' then
              \state\ <= get_wait2344;
            else
              \$602\ := \$603\;
              \$v2343\ := \$arr1451_ptr_take\;
              if \$v2343\(0) = '1' then
                \state\ <= q_wait2342;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$602\));
                \state\ <= pause_getI2340;
              end if;
            end if;
          when pause_getII2351 =>
            \$arr1452_ptr_take\(0) := '0';
            \$604\ := \$arr1452_value\;
            if \$604_lock\(0) = '1' then
              \state\ <= get_wait2349;
            else
              \$588\ := \$604\;
              \$v2348\ := \$arr1452_ptr_take\;
              if \$v2348\(0) = '1' then
                \state\ <= q_wait2347;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2345;
              end if;
            end if;
          when pause_getII2359 =>
            \$arr1451_ptr_take\(0) := '0';
            \$620\ := \$arr1451_value\;
            \$618\ := \$620\(36 to 71);
            \$v2356\ := \$618\;
            \$v2357\ := \$v2356\(0 to 3);
            \$v2355\ := \$v2356\(4 to 35);
            case \$v2357\ is
            when "0010" =>
              \$587\ := eclat_true;
              \$v2354\ := \$587\;
              if \$v2354\(0) = '1' then
                \$v2325\ := \$arr1452_ptr_take\;
                if \$v2325\(0) = '1' then
                  \state\ <= q_wait2324;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2322;
                end if;
              else
                \$v2353\ := \$arr1452_ptr_take\;
                if \$v2353\(0) = '1' then
                  \state\ <= q_wait2352;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2350;
                end if;
              end if;
            when others =>
              \$587\ := eclat_false;
              \$v2354\ := \$587\;
              if \$v2354\(0) = '1' then
                \$v2325\ := \$arr1452_ptr_take\;
                if \$v2325\(0) = '1' then
                  \state\ <= q_wait2324;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2322;
                end if;
              else
                \$v2353\ := \$arr1452_ptr_take\;
                if \$v2353\(0) = '1' then
                  \state\ <= q_wait2352;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2350;
                end if;
              end if;
            end case;
          when pause_getII2364 =>
            \$arr1452_ptr_take\(0) := '0';
            \$625\ := \$arr1452_value\;
            if \$625_lock\(0) = '1' then
              \state\ <= get_wait2362;
            else
              \$624\ := \$625\;
              \$v2361\ := \$arr1451_ptr_take\;
              if \$v2361\(0) = '1' then
                \state\ <= q_wait2360;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$624\));
                \state\ <= pause_getI2358;
              end if;
            end if;
          when pause_getII2368 =>
            \$arr1451_ptr_take\(0) := '0';
            \$626\ := \$arr1451_value\;
            \$586_x\ := \$626\(0 to 35);
            \$v2366\ := \$arr1452_ptr_take\;
            if \$v2366\(0) = '1' then
              \state\ <= q_wait2365;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2363;
            end if;
          when pause_getII2373 =>
            \$arr1452_ptr_take\(0) := '0';
            \$631\ := \$arr1452_value\;
            if \$631_lock\(0) = '1' then
              \state\ <= get_wait2371;
            else
              \$630\ := \$631\;
              \$v2370\ := \$arr1451_ptr_take\;
              if \$v2370\(0) = '1' then
                \state\ <= q_wait2369;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$630\));
                \state\ <= pause_getI2367;
              end if;
            end if;
          when pause_getII2383 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$640_lock\(0) = '1' then
              \state\ <= get_wait2380;
            else
              \$640_lock\ := eclat_true;
              \state\ <= get_pause2381;
            end if;
          when pause_getII2399 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$639_lock\(0) = '1' then
              \state\ <= get_wait2396;
            else
              \$639_lock\ := eclat_true;
              \state\ <= get_pause2397;
            end if;
          when pause_getII2422 =>
            \$arr1452_ptr_take\(0) := '0';
            \$641\ := \$arr1452_value\;
            if \$641_lock\(0) = '1' then
              \state\ <= get_wait2420;
            else
              \$635_i\ := \$641\;
              \$v2419\ := eclat_gt(\$635_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2419\(0) = '1' then
                \$v2418\ := eclat_eq(\$635_i\ & X"000" & X"15f90");
                if \$v2418\(0) = '1' then
                  \$v2395\ := \$arr1451_ptr_take\;
                  if \$v2395\(0) = '1' then
                    \state\ <= q_wait2394;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2389\ := "00000000000000000000000000000000";
                    \$v2390\ := "00000000000000000000000000000000";
                    \$v2391\ := "00000000000000000000000000000101";
                    \$v2386\ := "00000000000000000000000000000000";
                    \$v2387\ := "00000000000000000000000000000000";
                    \$v2388\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2389\ & "0001" & \$v2390\ & "0001" & \$v2391\ & "0001" & \$v2386\ & "0001" & \$v2387\ & "0001" & \$v2388\);
                    \state\ <= pause_setI2392;
                  end if;
                else
                  \$v2417\ := \$arr1451_ptr_take\;
                  if \$v2417\(0) = '1' then
                    \state\ <= q_wait2416;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v2411\ := "00000000000000000000000000000000";
                    \$v2412\ := "00000000000000000000000000000000";
                    \$v2413\ := "00000000000000000000000000000101";
                    \$v2408\ := "00000000000000000000000000000000";
                    \$v2409\ := "00000000000000000000000000000000";
                    \$v2410\ := "00000000000000000000000000000101";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2411\ & "0001" & \$v2412\ & "0001" & \$v2413\ & "0001" & \$v2408\ & "0001" & \$v2409\ & "0001" & \$v2410\);
                    \state\ <= pause_setI2414;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811413\;
              end if;
            end if;
          when pause_getII2440 =>
            \$arr1451_ptr_take\(0) := '0';
            \$668\ := \$arr1451_value\;
            \$663\ := \$668\(36 to 71);
            \$v2437\ := \$663\;
            \$v2438\ := \$v2437\(0 to 3);
            \$v2436\ := \$v2437\(4 to 35);
            case \$v2438\ is
            when "0010" =>
              \$664_i\ := \$v2436\(0 to 31);
              \$662\ := \$664_i\;
              if \$661_lock\(0) = '1' then
                \state\ <= get_wait2434;
              else
                \$661_lock\ := eclat_true;
                \state\ <= get_pause2435;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811414\;
            end case;
          when pause_getII2445 =>
            \$arr1452_ptr_take\(0) := '0';
            \$673\ := \$arr1452_value\;
            if \$673_lock\(0) = '1' then
              \state\ <= get_wait2443;
            else
              \$672\ := \$673\;
              \$v2442\ := \$arr1451_ptr_take\;
              if \$v2442\(0) = '1' then
                \state\ <= q_wait2441;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$672\));
                \state\ <= pause_getI2439;
              end if;
            end if;
          when pause_getII2449 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2447\ := \$arr1452_ptr_take\;
            if \$v2447\(0) = '1' then
              \state\ <= q_wait2446;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2444;
            end if;
          when pause_getII2458 =>
            \$arr1451_ptr_take\(0) := '0';
            \$648\ := \$arr1451_value\;
            \$647\ := \$648\(72 to 107);
            \$v2456\ := "00000000000000000000000000000000";
            \$645\ := "0000" & \$v2456\ & \$646\ & \$647\;
            \$v2455\ := \$arr1451_ptr_take\;
            if \$v2455\(0) = '1' then
              \state\ <= q_wait2454;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$644\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$645\;
              \state\ <= pause_setI2452;
            end if;
          when pause_getII2463 =>
            \$arr1452_ptr_take\(0) := '0';
            \$653\ := \$arr1452_value\;
            if \$653_lock\(0) = '1' then
              \state\ <= get_wait2461;
            else
              \$652\ := \$653\;
              \$v2460\ := \$arr1451_ptr_take\;
              if \$v2460\(0) = '1' then
                \state\ <= q_wait2459;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$652\));
                \state\ <= pause_getI2457;
              end if;
            end if;
          when pause_getII2467 =>
            \$arr1451_ptr_take\(0) := '0';
            \$654\ := \$arr1451_value\;
            \$646\ := \$654\(36 to 71);
            \$v2465\ := \$arr1452_ptr_take\;
            if \$v2465\(0) = '1' then
              \state\ <= q_wait2464;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2462;
            end if;
          when pause_getII2472 =>
            \$arr1452_ptr_take\(0) := '0';
            \$659\ := \$arr1452_value\;
            if \$659_lock\(0) = '1' then
              \state\ <= get_wait2470;
            else
              \$658\ := \$659\;
              \$v2469\ := \$arr1451_ptr_take\;
              if \$v2469\(0) = '1' then
                \state\ <= q_wait2468;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$658\));
                \state\ <= pause_getI2466;
              end if;
            end if;
          when pause_getII2477 =>
            \$arr1452_ptr_take\(0) := '0';
            \$660\ := \$arr1452_value\;
            if \$660_lock\(0) = '1' then
              \state\ <= get_wait2475;
            else
              \$644\ := \$660\;
              \$v2474\ := \$arr1452_ptr_take\;
              if \$v2474\(0) = '1' then
                \state\ <= q_wait2473;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2471;
              end if;
            end if;
          when pause_getII2485 =>
            \$arr1451_ptr_take\(0) := '0';
            \$676\ := \$arr1451_value\;
            \$674\ := \$676\(36 to 71);
            \$v2482\ := \$674\;
            \$v2483\ := \$v2482\(0 to 3);
            \$v2481\ := \$v2482\(4 to 35);
            case \$v2483\ is
            when "0010" =>
              \$643\ := eclat_true;
              \$v2480\ := \$643\;
              if \$v2480\(0) = '1' then
                \$v2451\ := \$arr1452_ptr_take\;
                if \$v2451\(0) = '1' then
                  \state\ <= q_wait2450;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2448;
                end if;
              else
                \$v2479\ := \$arr1452_ptr_take\;
                if \$v2479\(0) = '1' then
                  \state\ <= q_wait2478;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2476;
                end if;
              end if;
            when others =>
              \$643\ := eclat_false;
              \$v2480\ := \$643\;
              if \$v2480\(0) = '1' then
                \$v2451\ := \$arr1452_ptr_take\;
                if \$v2451\(0) = '1' then
                  \state\ <= q_wait2450;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2448;
                end if;
              else
                \$v2479\ := \$arr1452_ptr_take\;
                if \$v2479\(0) = '1' then
                  \state\ <= q_wait2478;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2476;
                end if;
              end if;
            end case;
          when pause_getII2490 =>
            \$arr1452_ptr_take\(0) := '0';
            \$681\ := \$arr1452_value\;
            if \$681_lock\(0) = '1' then
              \state\ <= get_wait2488;
            else
              \$680\ := \$681\;
              \$v2487\ := \$arr1451_ptr_take\;
              if \$v2487\(0) = '1' then
                \state\ <= q_wait2486;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$680\));
                \state\ <= pause_getI2484;
              end if;
            end if;
          when pause_getII2494 =>
            \$arr1451_ptr_take\(0) := '0';
            \$682\ := \$arr1451_value\;
            \$642_x\ := \$682\(0 to 35);
            \$v2492\ := \$arr1452_ptr_take\;
            if \$v2492\(0) = '1' then
              \state\ <= q_wait2491;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2489;
            end if;
          when pause_getII2499 =>
            \$arr1452_ptr_take\(0) := '0';
            \$687\ := \$arr1452_value\;
            if \$687_lock\(0) = '1' then
              \state\ <= get_wait2497;
            else
              \$686\ := \$687\;
              \$v2496\ := \$arr1451_ptr_take\;
              if \$v2496\(0) = '1' then
                \state\ <= q_wait2495;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$686\));
                \state\ <= pause_getI2493;
              end if;
            end if;
          when pause_getII2508 =>
            \$arr1451_ptr_take\(0) := '0';
            \$714\ := \$arr1451_value\;
            \$709\ := \$714\(36 to 71);
            \$v2505\ := \$709\;
            \$v2506\ := \$v2505\(0 to 3);
            \$v2504\ := \$v2505\(4 to 35);
            case \$v2506\ is
            when "0010" =>
              \$710_i\ := \$v2504\(0 to 31);
              \$708\ := \$710_i\;
              if \$707_lock\(0) = '1' then
                \state\ <= get_wait2502;
              else
                \$707_lock\ := eclat_true;
                \state\ <= get_pause2503;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811415\;
            end case;
          when pause_getII2513 =>
            \$arr1452_ptr_take\(0) := '0';
            \$719\ := \$arr1452_value\;
            if \$719_lock\(0) = '1' then
              \state\ <= get_wait2511;
            else
              \$718\ := \$719\;
              \$v2510\ := \$arr1451_ptr_take\;
              if \$v2510\(0) = '1' then
                \state\ <= q_wait2509;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$718\));
                \state\ <= pause_getI2507;
              end if;
            end if;
          when pause_getII2517 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2515\ := \$arr1452_ptr_take\;
            if \$v2515\(0) = '1' then
              \state\ <= q_wait2514;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2512;
            end if;
          when pause_getII2526 =>
            \$arr1451_ptr_take\(0) := '0';
            \$694\ := \$arr1451_value\;
            \$693\ := \$694\(72 to 107);
            \$v2524\ := "00000000000000000000000000000000";
            \$691\ := "0000" & \$v2524\ & \$692\ & \$693\;
            \$v2523\ := \$arr1451_ptr_take\;
            if \$v2523\(0) = '1' then
              \state\ <= q_wait2522;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$690\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$691\;
              \state\ <= pause_setI2520;
            end if;
          when pause_getII2531 =>
            \$arr1452_ptr_take\(0) := '0';
            \$699\ := \$arr1452_value\;
            if \$699_lock\(0) = '1' then
              \state\ <= get_wait2529;
            else
              \$698\ := \$699\;
              \$v2528\ := \$arr1451_ptr_take\;
              if \$v2528\(0) = '1' then
                \state\ <= q_wait2527;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$698\));
                \state\ <= pause_getI2525;
              end if;
            end if;
          when pause_getII2535 =>
            \$arr1451_ptr_take\(0) := '0';
            \$700\ := \$arr1451_value\;
            \$692\ := \$700\(36 to 71);
            \$v2533\ := \$arr1452_ptr_take\;
            if \$v2533\(0) = '1' then
              \state\ <= q_wait2532;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2530;
            end if;
          when pause_getII2540 =>
            \$arr1452_ptr_take\(0) := '0';
            \$705\ := \$arr1452_value\;
            if \$705_lock\(0) = '1' then
              \state\ <= get_wait2538;
            else
              \$704\ := \$705\;
              \$v2537\ := \$arr1451_ptr_take\;
              if \$v2537\(0) = '1' then
                \state\ <= q_wait2536;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$704\));
                \state\ <= pause_getI2534;
              end if;
            end if;
          when pause_getII2545 =>
            \$arr1452_ptr_take\(0) := '0';
            \$706\ := \$arr1452_value\;
            if \$706_lock\(0) = '1' then
              \state\ <= get_wait2543;
            else
              \$690\ := \$706\;
              \$v2542\ := \$arr1452_ptr_take\;
              if \$v2542\(0) = '1' then
                \state\ <= q_wait2541;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2539;
              end if;
            end if;
          when pause_getII2553 =>
            \$arr1451_ptr_take\(0) := '0';
            \$722\ := \$arr1451_value\;
            \$720\ := \$722\(36 to 71);
            \$v2550\ := \$720\;
            \$v2551\ := \$v2550\(0 to 3);
            \$v2549\ := \$v2550\(4 to 35);
            case \$v2551\ is
            when "0010" =>
              \$689\ := eclat_true;
              \$v2548\ := \$689\;
              if \$v2548\(0) = '1' then
                \$v2519\ := \$arr1452_ptr_take\;
                if \$v2519\(0) = '1' then
                  \state\ <= q_wait2518;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2516;
                end if;
              else
                \$v2547\ := \$arr1452_ptr_take\;
                if \$v2547\(0) = '1' then
                  \state\ <= q_wait2546;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2544;
                end if;
              end if;
            when others =>
              \$689\ := eclat_false;
              \$v2548\ := \$689\;
              if \$v2548\(0) = '1' then
                \$v2519\ := \$arr1452_ptr_take\;
                if \$v2519\(0) = '1' then
                  \state\ <= q_wait2518;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2516;
                end if;
              else
                \$v2547\ := \$arr1452_ptr_take\;
                if \$v2547\(0) = '1' then
                  \state\ <= q_wait2546;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2544;
                end if;
              end if;
            end case;
          when pause_getII2558 =>
            \$arr1452_ptr_take\(0) := '0';
            \$727\ := \$arr1452_value\;
            if \$727_lock\(0) = '1' then
              \state\ <= get_wait2556;
            else
              \$726\ := \$727\;
              \$v2555\ := \$arr1451_ptr_take\;
              if \$v2555\(0) = '1' then
                \state\ <= q_wait2554;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$726\));
                \state\ <= pause_getI2552;
              end if;
            end if;
          when pause_getII2562 =>
            \$arr1451_ptr_take\(0) := '0';
            \$728\ := \$arr1451_value\;
            \$688_x\ := \$728\(0 to 35);
            \$v2560\ := \$arr1452_ptr_take\;
            if \$v2560\(0) = '1' then
              \state\ <= q_wait2559;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2557;
            end if;
          when pause_getII2567 =>
            \$arr1452_ptr_take\(0) := '0';
            \$733\ := \$arr1452_value\;
            if \$733_lock\(0) = '1' then
              \state\ <= get_wait2565;
            else
              \$732\ := \$733\;
              \$v2564\ := \$arr1451_ptr_take\;
              if \$v2564\(0) = '1' then
                \state\ <= q_wait2563;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$732\));
                \state\ <= pause_getI2561;
              end if;
            end if;
          when pause_getII2577 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$739_lock\(0) = '1' then
              \state\ <= get_wait2574;
            else
              \$739_lock\ := eclat_true;
              \state\ <= get_pause2575;
            end if;
          when pause_getII2587 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$738_lock\(0) = '1' then
              \state\ <= get_wait2584;
            else
              \$738_lock\ := eclat_true;
              \state\ <= get_pause2585;
            end if;
          when pause_getII2604 =>
            \$arr1452_ptr_take\(0) := '0';
            \$743\ := \$arr1452_value\;
            if \$743_lock\(0) = '1' then
              \state\ <= get_wait2602;
            else
              \$734_i\ := \$743\;
              \$v2601\ := eclat_gt(\$734_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2601\(0) = '1' then
                \$v2600\ := eclat_eq(\$734_i\ & X"000" & X"15f90");
                if \$v2600\(0) = '1' then
                  \$v2583\ := \$arr1451_ptr_take\;
                  if \$v2583\(0) = '1' then
                    \state\ <= q_wait2582;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
                    \state\ <= pause_setI2580;
                  end if;
                else
                  \$v2599\ := \$arr1451_ptr_take\;
                  if \$v2599\(0) = '1' then
                    \state\ <= q_wait2598;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
                    \state\ <= pause_setI2596;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811416\;
              end if;
            end if;
          when pause_getII2609 =>
            \$arr1451_ptr_take\(0) := '0';
            \$56_y\ := \$arr1451_value\;
            \$v2606\ := \$arr1452_ptr_take\;
            if \$v2606\(0) = '1' then
              \state\ <= q_wait2605;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2603;
            end if;
          when pause_getII2620 =>
            \$arr1451_ptr_take\(0) := '0';
            \$773\ := \$arr1451_value\;
            \$768\ := \$773\(36 to 71);
            \$v2617\ := \$768\;
            \$v2618\ := \$v2617\(0 to 3);
            \$v2616\ := \$v2617\(4 to 35);
            case \$v2618\ is
            when "0010" =>
              \$769_i\ := \$v2616\(0 to 31);
              \$767\ := \$769_i\;
              if \$766_lock\(0) = '1' then
                \state\ <= get_wait2614;
              else
                \$766_lock\ := eclat_true;
                \state\ <= get_pause2615;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811418\;
            end case;
          when pause_getII2625 =>
            \$arr1452_ptr_take\(0) := '0';
            \$778\ := \$arr1452_value\;
            if \$778_lock\(0) = '1' then
              \state\ <= get_wait2623;
            else
              \$777\ := \$778\;
              \$v2622\ := \$arr1451_ptr_take\;
              if \$v2622\(0) = '1' then
                \state\ <= q_wait2621;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$777\));
                \state\ <= pause_getI2619;
              end if;
            end if;
          when pause_getII2629 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2627\ := \$arr1452_ptr_take\;
            if \$v2627\(0) = '1' then
              \state\ <= q_wait2626;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2624;
            end if;
          when pause_getII2638 =>
            \$arr1451_ptr_take\(0) := '0';
            \$753\ := \$arr1451_value\;
            \$752\ := \$753\(72 to 107);
            \$v2636\ := "00000000000000000000000000000000";
            \$750\ := "0000" & \$v2636\ & \$751\ & \$752\;
            \$v2635\ := \$arr1451_ptr_take\;
            if \$v2635\(0) = '1' then
              \state\ <= q_wait2634;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$749\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$750\;
              \state\ <= pause_setI2632;
            end if;
          when pause_getII2643 =>
            \$arr1452_ptr_take\(0) := '0';
            \$758\ := \$arr1452_value\;
            if \$758_lock\(0) = '1' then
              \state\ <= get_wait2641;
            else
              \$757\ := \$758\;
              \$v2640\ := \$arr1451_ptr_take\;
              if \$v2640\(0) = '1' then
                \state\ <= q_wait2639;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$757\));
                \state\ <= pause_getI2637;
              end if;
            end if;
          when pause_getII2647 =>
            \$arr1451_ptr_take\(0) := '0';
            \$759\ := \$arr1451_value\;
            \$751\ := \$759\(36 to 71);
            \$v2645\ := \$arr1452_ptr_take\;
            if \$v2645\(0) = '1' then
              \state\ <= q_wait2644;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2642;
            end if;
          when pause_getII2652 =>
            \$arr1452_ptr_take\(0) := '0';
            \$764\ := \$arr1452_value\;
            if \$764_lock\(0) = '1' then
              \state\ <= get_wait2650;
            else
              \$763\ := \$764\;
              \$v2649\ := \$arr1451_ptr_take\;
              if \$v2649\(0) = '1' then
                \state\ <= q_wait2648;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$763\));
                \state\ <= pause_getI2646;
              end if;
            end if;
          when pause_getII2657 =>
            \$arr1452_ptr_take\(0) := '0';
            \$765\ := \$arr1452_value\;
            if \$765_lock\(0) = '1' then
              \state\ <= get_wait2655;
            else
              \$749\ := \$765\;
              \$v2654\ := \$arr1452_ptr_take\;
              if \$v2654\(0) = '1' then
                \state\ <= q_wait2653;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2651;
              end if;
            end if;
          when pause_getII2665 =>
            \$arr1451_ptr_take\(0) := '0';
            \$781\ := \$arr1451_value\;
            \$779\ := \$781\(36 to 71);
            \$v2662\ := \$779\;
            \$v2663\ := \$v2662\(0 to 3);
            \$v2661\ := \$v2662\(4 to 35);
            case \$v2663\ is
            when "0010" =>
              \$748\ := eclat_true;
              \$v2660\ := \$748\;
              if \$v2660\(0) = '1' then
                \$v2631\ := \$arr1452_ptr_take\;
                if \$v2631\(0) = '1' then
                  \state\ <= q_wait2630;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2628;
                end if;
              else
                \$v2659\ := \$arr1452_ptr_take\;
                if \$v2659\(0) = '1' then
                  \state\ <= q_wait2658;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2656;
                end if;
              end if;
            when others =>
              \$748\ := eclat_false;
              \$v2660\ := \$748\;
              if \$v2660\(0) = '1' then
                \$v2631\ := \$arr1452_ptr_take\;
                if \$v2631\(0) = '1' then
                  \state\ <= q_wait2630;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2628;
                end if;
              else
                \$v2659\ := \$arr1452_ptr_take\;
                if \$v2659\(0) = '1' then
                  \state\ <= q_wait2658;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2656;
                end if;
              end if;
            end case;
          when pause_getII2670 =>
            \$arr1452_ptr_take\(0) := '0';
            \$786\ := \$arr1452_value\;
            if \$786_lock\(0) = '1' then
              \state\ <= get_wait2668;
            else
              \$785\ := \$786\;
              \$v2667\ := \$arr1451_ptr_take\;
              if \$v2667\(0) = '1' then
                \state\ <= q_wait2666;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$785\));
                \state\ <= pause_getI2664;
              end if;
            end if;
          when pause_getII2674 =>
            \$arr1451_ptr_take\(0) := '0';
            \$787\ := \$arr1451_value\;
            \$747_x\ := \$787\(0 to 35);
            \$v2672\ := \$arr1452_ptr_take\;
            if \$v2672\(0) = '1' then
              \state\ <= q_wait2671;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2669;
            end if;
          when pause_getII2679 =>
            \$arr1452_ptr_take\(0) := '0';
            \$792\ := \$arr1452_value\;
            if \$792_lock\(0) = '1' then
              \state\ <= get_wait2677;
            else
              \$791\ := \$792\;
              \$v2676\ := \$arr1451_ptr_take\;
              if \$v2676\(0) = '1' then
                \state\ <= q_wait2675;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$791\));
                \state\ <= pause_getI2673;
              end if;
            end if;
          when pause_getII2688 =>
            \$arr1451_ptr_take\(0) := '0';
            \$819\ := \$arr1451_value\;
            \$814\ := \$819\(36 to 71);
            \$v2685\ := \$814\;
            \$v2686\ := \$v2685\(0 to 3);
            \$v2684\ := \$v2685\(4 to 35);
            case \$v2686\ is
            when "0010" =>
              \$815_i\ := \$v2684\(0 to 31);
              \$813\ := \$815_i\;
              if \$812_lock\(0) = '1' then
                \state\ <= get_wait2682;
              else
                \$812_lock\ := eclat_true;
                \state\ <= get_pause2683;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811419\;
            end case;
          when pause_getII2693 =>
            \$arr1452_ptr_take\(0) := '0';
            \$824\ := \$arr1452_value\;
            if \$824_lock\(0) = '1' then
              \state\ <= get_wait2691;
            else
              \$823\ := \$824\;
              \$v2690\ := \$arr1451_ptr_take\;
              if \$v2690\(0) = '1' then
                \state\ <= q_wait2689;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$823\));
                \state\ <= pause_getI2687;
              end if;
            end if;
          when pause_getII2697 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2695\ := \$arr1452_ptr_take\;
            if \$v2695\(0) = '1' then
              \state\ <= q_wait2694;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2692;
            end if;
          when pause_getII2706 =>
            \$arr1451_ptr_take\(0) := '0';
            \$799\ := \$arr1451_value\;
            \$798\ := \$799\(72 to 107);
            \$v2704\ := "00000000000000000000000000000000";
            \$796\ := "0000" & \$v2704\ & \$797\ & \$798\;
            \$v2703\ := \$arr1451_ptr_take\;
            if \$v2703\(0) = '1' then
              \state\ <= q_wait2702;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$795\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$796\;
              \state\ <= pause_setI2700;
            end if;
          when pause_getII2711 =>
            \$arr1452_ptr_take\(0) := '0';
            \$804\ := \$arr1452_value\;
            if \$804_lock\(0) = '1' then
              \state\ <= get_wait2709;
            else
              \$803\ := \$804\;
              \$v2708\ := \$arr1451_ptr_take\;
              if \$v2708\(0) = '1' then
                \state\ <= q_wait2707;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$803\));
                \state\ <= pause_getI2705;
              end if;
            end if;
          when pause_getII2715 =>
            \$arr1451_ptr_take\(0) := '0';
            \$805\ := \$arr1451_value\;
            \$797\ := \$805\(36 to 71);
            \$v2713\ := \$arr1452_ptr_take\;
            if \$v2713\(0) = '1' then
              \state\ <= q_wait2712;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2710;
            end if;
          when pause_getII2720 =>
            \$arr1452_ptr_take\(0) := '0';
            \$810\ := \$arr1452_value\;
            if \$810_lock\(0) = '1' then
              \state\ <= get_wait2718;
            else
              \$809\ := \$810\;
              \$v2717\ := \$arr1451_ptr_take\;
              if \$v2717\(0) = '1' then
                \state\ <= q_wait2716;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$809\));
                \state\ <= pause_getI2714;
              end if;
            end if;
          when pause_getII2725 =>
            \$arr1452_ptr_take\(0) := '0';
            \$811\ := \$arr1452_value\;
            if \$811_lock\(0) = '1' then
              \state\ <= get_wait2723;
            else
              \$795\ := \$811\;
              \$v2722\ := \$arr1452_ptr_take\;
              if \$v2722\(0) = '1' then
                \state\ <= q_wait2721;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2719;
              end if;
            end if;
          when pause_getII2733 =>
            \$arr1451_ptr_take\(0) := '0';
            \$827\ := \$arr1451_value\;
            \$825\ := \$827\(36 to 71);
            \$v2730\ := \$825\;
            \$v2731\ := \$v2730\(0 to 3);
            \$v2729\ := \$v2730\(4 to 35);
            case \$v2731\ is
            when "0010" =>
              \$794\ := eclat_true;
              \$v2728\ := \$794\;
              if \$v2728\(0) = '1' then
                \$v2699\ := \$arr1452_ptr_take\;
                if \$v2699\(0) = '1' then
                  \state\ <= q_wait2698;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2696;
                end if;
              else
                \$v2727\ := \$arr1452_ptr_take\;
                if \$v2727\(0) = '1' then
                  \state\ <= q_wait2726;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2724;
                end if;
              end if;
            when others =>
              \$794\ := eclat_false;
              \$v2728\ := \$794\;
              if \$v2728\(0) = '1' then
                \$v2699\ := \$arr1452_ptr_take\;
                if \$v2699\(0) = '1' then
                  \state\ <= q_wait2698;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2696;
                end if;
              else
                \$v2727\ := \$arr1452_ptr_take\;
                if \$v2727\(0) = '1' then
                  \state\ <= q_wait2726;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2724;
                end if;
              end if;
            end case;
          when pause_getII2738 =>
            \$arr1452_ptr_take\(0) := '0';
            \$832\ := \$arr1452_value\;
            if \$832_lock\(0) = '1' then
              \state\ <= get_wait2736;
            else
              \$831\ := \$832\;
              \$v2735\ := \$arr1451_ptr_take\;
              if \$v2735\(0) = '1' then
                \state\ <= q_wait2734;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$831\));
                \state\ <= pause_getI2732;
              end if;
            end if;
          when pause_getII2742 =>
            \$arr1451_ptr_take\(0) := '0';
            \$833\ := \$arr1451_value\;
            \$793_x\ := \$833\(0 to 35);
            \$v2740\ := \$arr1452_ptr_take\;
            if \$v2740\(0) = '1' then
              \state\ <= q_wait2739;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2737;
            end if;
          when pause_getII2747 =>
            \$arr1452_ptr_take\(0) := '0';
            \$838\ := \$arr1452_value\;
            if \$838_lock\(0) = '1' then
              \state\ <= get_wait2745;
            else
              \$837\ := \$838\;
              \$v2744\ := \$arr1451_ptr_take\;
              if \$v2744\(0) = '1' then
                \state\ <= q_wait2743;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$837\));
                \state\ <= pause_getI2741;
              end if;
            end if;
          when pause_getII2757 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$846_lock\(0) = '1' then
              \state\ <= get_wait2754;
            else
              \$846_lock\ := eclat_true;
              \state\ <= get_pause2755;
            end if;
          when pause_getII2767 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$845_lock\(0) = '1' then
              \state\ <= get_wait2764;
            else
              \$845_lock\ := eclat_true;
              \state\ <= get_pause2765;
            end if;
          when pause_getII2784 =>
            \$arr1452_ptr_take\(0) := '0';
            \$850\ := \$arr1452_value\;
            if \$850_lock\(0) = '1' then
              \state\ <= get_wait2782;
            else
              \$841_i\ := \$850\;
              \$v2781\ := eclat_gt(\$841_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2781\(0) = '1' then
                \$v2780\ := eclat_eq(\$841_i\ & X"000" & X"15f90");
                if \$v2780\(0) = '1' then
                  \$v2763\ := \$arr1451_ptr_take\;
                  if \$v2763\(0) = '1' then
                    \state\ <= q_wait2762;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
                    \state\ <= pause_setI2760;
                  end if;
                else
                  \$v2779\ := \$arr1451_ptr_take\;
                  if \$v2779\(0) = '1' then
                    \state\ <= q_wait2778;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
                    \state\ <= pause_setI2776;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811420\;
              end if;
            end if;
          when pause_getII2789 =>
            \$arr1451_ptr_take\(0) := '0';
            \$840_y\ := \$arr1451_value\;
            \$v2786\ := \$arr1452_ptr_take\;
            if \$v2786\(0) = '1' then
              \state\ <= q_wait2785;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2783;
            end if;
          when pause_getII2800 =>
            \$arr1451_ptr_take\(0) := '0';
            \$882\ := \$arr1451_value\;
            \$877\ := \$882\(36 to 71);
            \$v2797\ := \$877\;
            \$v2798\ := \$v2797\(0 to 3);
            \$v2796\ := \$v2797\(4 to 35);
            case \$v2798\ is
            when "0010" =>
              \$878_i\ := \$v2796\(0 to 31);
              \$876\ := \$878_i\;
              if \$875_lock\(0) = '1' then
                \state\ <= get_wait2794;
              else
                \$875_lock\ := eclat_true;
                \state\ <= get_pause2795;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811422\;
            end case;
          when pause_getII2805 =>
            \$arr1452_ptr_take\(0) := '0';
            \$887\ := \$arr1452_value\;
            if \$887_lock\(0) = '1' then
              \state\ <= get_wait2803;
            else
              \$886\ := \$887\;
              \$v2802\ := \$arr1451_ptr_take\;
              if \$v2802\(0) = '1' then
                \state\ <= q_wait2801;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$886\));
                \state\ <= pause_getI2799;
              end if;
            end if;
          when pause_getII2809 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2807\ := \$arr1452_ptr_take\;
            if \$v2807\(0) = '1' then
              \state\ <= q_wait2806;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2804;
            end if;
          when pause_getII2818 =>
            \$arr1451_ptr_take\(0) := '0';
            \$862\ := \$arr1451_value\;
            \$861\ := \$862\(72 to 107);
            \$v2816\ := "00000000000000000000000000000000";
            \$859\ := "0000" & \$v2816\ & \$860\ & \$861\;
            \$v2815\ := \$arr1451_ptr_take\;
            if \$v2815\(0) = '1' then
              \state\ <= q_wait2814;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$858\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$859\;
              \state\ <= pause_setI2812;
            end if;
          when pause_getII2823 =>
            \$arr1452_ptr_take\(0) := '0';
            \$867\ := \$arr1452_value\;
            if \$867_lock\(0) = '1' then
              \state\ <= get_wait2821;
            else
              \$866\ := \$867\;
              \$v2820\ := \$arr1451_ptr_take\;
              if \$v2820\(0) = '1' then
                \state\ <= q_wait2819;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$866\));
                \state\ <= pause_getI2817;
              end if;
            end if;
          when pause_getII2827 =>
            \$arr1451_ptr_take\(0) := '0';
            \$868\ := \$arr1451_value\;
            \$860\ := \$868\(36 to 71);
            \$v2825\ := \$arr1452_ptr_take\;
            if \$v2825\(0) = '1' then
              \state\ <= q_wait2824;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2822;
            end if;
          when pause_getII2832 =>
            \$arr1452_ptr_take\(0) := '0';
            \$873\ := \$arr1452_value\;
            if \$873_lock\(0) = '1' then
              \state\ <= get_wait2830;
            else
              \$872\ := \$873\;
              \$v2829\ := \$arr1451_ptr_take\;
              if \$v2829\(0) = '1' then
                \state\ <= q_wait2828;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$872\));
                \state\ <= pause_getI2826;
              end if;
            end if;
          when pause_getII2837 =>
            \$arr1452_ptr_take\(0) := '0';
            \$874\ := \$arr1452_value\;
            if \$874_lock\(0) = '1' then
              \state\ <= get_wait2835;
            else
              \$858\ := \$874\;
              \$v2834\ := \$arr1452_ptr_take\;
              if \$v2834\(0) = '1' then
                \state\ <= q_wait2833;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2831;
              end if;
            end if;
          when pause_getII2845 =>
            \$arr1451_ptr_take\(0) := '0';
            \$890\ := \$arr1451_value\;
            \$888\ := \$890\(36 to 71);
            \$v2842\ := \$888\;
            \$v2843\ := \$v2842\(0 to 3);
            \$v2841\ := \$v2842\(4 to 35);
            case \$v2843\ is
            when "0010" =>
              \$857\ := eclat_true;
              \$v2840\ := \$857\;
              if \$v2840\(0) = '1' then
                \$v2811\ := \$arr1452_ptr_take\;
                if \$v2811\(0) = '1' then
                  \state\ <= q_wait2810;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2808;
                end if;
              else
                \$v2839\ := \$arr1452_ptr_take\;
                if \$v2839\(0) = '1' then
                  \state\ <= q_wait2838;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2836;
                end if;
              end if;
            when others =>
              \$857\ := eclat_false;
              \$v2840\ := \$857\;
              if \$v2840\(0) = '1' then
                \$v2811\ := \$arr1452_ptr_take\;
                if \$v2811\(0) = '1' then
                  \state\ <= q_wait2810;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2808;
                end if;
              else
                \$v2839\ := \$arr1452_ptr_take\;
                if \$v2839\(0) = '1' then
                  \state\ <= q_wait2838;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2836;
                end if;
              end if;
            end case;
          when pause_getII2850 =>
            \$arr1452_ptr_take\(0) := '0';
            \$895\ := \$arr1452_value\;
            if \$895_lock\(0) = '1' then
              \state\ <= get_wait2848;
            else
              \$894\ := \$895\;
              \$v2847\ := \$arr1451_ptr_take\;
              if \$v2847\(0) = '1' then
                \state\ <= q_wait2846;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$894\));
                \state\ <= pause_getI2844;
              end if;
            end if;
          when pause_getII2854 =>
            \$arr1451_ptr_take\(0) := '0';
            \$896\ := \$arr1451_value\;
            \$856_x\ := \$896\(0 to 35);
            \$v2852\ := \$arr1452_ptr_take\;
            if \$v2852\(0) = '1' then
              \state\ <= q_wait2851;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2849;
            end if;
          when pause_getII2859 =>
            \$arr1452_ptr_take\(0) := '0';
            \$901\ := \$arr1452_value\;
            if \$901_lock\(0) = '1' then
              \state\ <= get_wait2857;
            else
              \$900\ := \$901\;
              \$v2856\ := \$arr1451_ptr_take\;
              if \$v2856\(0) = '1' then
                \state\ <= q_wait2855;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$900\));
                \state\ <= pause_getI2853;
              end if;
            end if;
          when pause_getII2868 =>
            \$arr1451_ptr_take\(0) := '0';
            \$928\ := \$arr1451_value\;
            \$923\ := \$928\(36 to 71);
            \$v2865\ := \$923\;
            \$v2866\ := \$v2865\(0 to 3);
            \$v2864\ := \$v2865\(4 to 35);
            case \$v2866\ is
            when "0010" =>
              \$924_i\ := \$v2864\(0 to 31);
              \$922\ := \$924_i\;
              if \$921_lock\(0) = '1' then
                \state\ <= get_wait2862;
              else
                \$921_lock\ := eclat_true;
                \state\ <= get_pause2863;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811423\;
            end case;
          when pause_getII2873 =>
            \$arr1452_ptr_take\(0) := '0';
            \$933\ := \$arr1452_value\;
            if \$933_lock\(0) = '1' then
              \state\ <= get_wait2871;
            else
              \$932\ := \$933\;
              \$v2870\ := \$arr1451_ptr_take\;
              if \$v2870\(0) = '1' then
                \state\ <= q_wait2869;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$932\));
                \state\ <= pause_getI2867;
              end if;
            end if;
          when pause_getII2877 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2875\ := \$arr1452_ptr_take\;
            if \$v2875\(0) = '1' then
              \state\ <= q_wait2874;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2872;
            end if;
          when pause_getII2886 =>
            \$arr1451_ptr_take\(0) := '0';
            \$908\ := \$arr1451_value\;
            \$907\ := \$908\(72 to 107);
            \$v2884\ := "00000000000000000000000000000000";
            \$905\ := "0000" & \$v2884\ & \$906\ & \$907\;
            \$v2883\ := \$arr1451_ptr_take\;
            if \$v2883\(0) = '1' then
              \state\ <= q_wait2882;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$904\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$905\;
              \state\ <= pause_setI2880;
            end if;
          when pause_getII2891 =>
            \$arr1452_ptr_take\(0) := '0';
            \$913\ := \$arr1452_value\;
            if \$913_lock\(0) = '1' then
              \state\ <= get_wait2889;
            else
              \$912\ := \$913\;
              \$v2888\ := \$arr1451_ptr_take\;
              if \$v2888\(0) = '1' then
                \state\ <= q_wait2887;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$912\));
                \state\ <= pause_getI2885;
              end if;
            end if;
          when pause_getII2895 =>
            \$arr1451_ptr_take\(0) := '0';
            \$914\ := \$arr1451_value\;
            \$906\ := \$914\(36 to 71);
            \$v2893\ := \$arr1452_ptr_take\;
            if \$v2893\(0) = '1' then
              \state\ <= q_wait2892;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2890;
            end if;
          when pause_getII2900 =>
            \$arr1452_ptr_take\(0) := '0';
            \$919\ := \$arr1452_value\;
            if \$919_lock\(0) = '1' then
              \state\ <= get_wait2898;
            else
              \$918\ := \$919\;
              \$v2897\ := \$arr1451_ptr_take\;
              if \$v2897\(0) = '1' then
                \state\ <= q_wait2896;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$918\));
                \state\ <= pause_getI2894;
              end if;
            end if;
          when pause_getII2905 =>
            \$arr1452_ptr_take\(0) := '0';
            \$920\ := \$arr1452_value\;
            if \$920_lock\(0) = '1' then
              \state\ <= get_wait2903;
            else
              \$904\ := \$920\;
              \$v2902\ := \$arr1452_ptr_take\;
              if \$v2902\(0) = '1' then
                \state\ <= q_wait2901;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2899;
              end if;
            end if;
          when pause_getII2913 =>
            \$arr1451_ptr_take\(0) := '0';
            \$936\ := \$arr1451_value\;
            \$934\ := \$936\(36 to 71);
            \$v2910\ := \$934\;
            \$v2911\ := \$v2910\(0 to 3);
            \$v2909\ := \$v2910\(4 to 35);
            case \$v2911\ is
            when "0010" =>
              \$903\ := eclat_true;
              \$v2908\ := \$903\;
              if \$v2908\(0) = '1' then
                \$v2879\ := \$arr1452_ptr_take\;
                if \$v2879\(0) = '1' then
                  \state\ <= q_wait2878;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2876;
                end if;
              else
                \$v2907\ := \$arr1452_ptr_take\;
                if \$v2907\(0) = '1' then
                  \state\ <= q_wait2906;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2904;
                end if;
              end if;
            when others =>
              \$903\ := eclat_false;
              \$v2908\ := \$903\;
              if \$v2908\(0) = '1' then
                \$v2879\ := \$arr1452_ptr_take\;
                if \$v2879\(0) = '1' then
                  \state\ <= q_wait2878;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2876;
                end if;
              else
                \$v2907\ := \$arr1452_ptr_take\;
                if \$v2907\(0) = '1' then
                  \state\ <= q_wait2906;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2904;
                end if;
              end if;
            end case;
          when pause_getII2918 =>
            \$arr1452_ptr_take\(0) := '0';
            \$941\ := \$arr1452_value\;
            if \$941_lock\(0) = '1' then
              \state\ <= get_wait2916;
            else
              \$940\ := \$941\;
              \$v2915\ := \$arr1451_ptr_take\;
              if \$v2915\(0) = '1' then
                \state\ <= q_wait2914;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$940\));
                \state\ <= pause_getI2912;
              end if;
            end if;
          when pause_getII2922 =>
            \$arr1451_ptr_take\(0) := '0';
            \$942\ := \$arr1451_value\;
            \$902_x\ := \$942\(0 to 35);
            \$v2920\ := \$arr1452_ptr_take\;
            if \$v2920\(0) = '1' then
              \state\ <= q_wait2919;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2917;
            end if;
          when pause_getII2927 =>
            \$arr1452_ptr_take\(0) := '0';
            \$947\ := \$arr1452_value\;
            if \$947_lock\(0) = '1' then
              \state\ <= get_wait2925;
            else
              \$946\ := \$947\;
              \$v2924\ := \$arr1451_ptr_take\;
              if \$v2924\(0) = '1' then
                \state\ <= q_wait2923;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$946\));
                \state\ <= pause_getI2921;
              end if;
            end if;
          when pause_getII2937 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$955_lock\(0) = '1' then
              \state\ <= get_wait2934;
            else
              \$955_lock\ := eclat_true;
              \state\ <= get_pause2935;
            end if;
          when pause_getII2947 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$954_lock\(0) = '1' then
              \state\ <= get_wait2944;
            else
              \$954_lock\ := eclat_true;
              \state\ <= get_pause2945;
            end if;
          when pause_getII2964 =>
            \$arr1452_ptr_take\(0) := '0';
            \$959\ := \$arr1452_value\;
            if \$959_lock\(0) = '1' then
              \state\ <= get_wait2962;
            else
              \$950_i\ := \$959\;
              \$v2961\ := eclat_gt(\$950_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v2961\(0) = '1' then
                \$v2960\ := eclat_eq(\$950_i\ & X"000" & X"15f90");
                if \$v2960\(0) = '1' then
                  \$v2943\ := \$arr1451_ptr_take\;
                  if \$v2943\(0) = '1' then
                    \state\ <= q_wait2942;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
                    \state\ <= pause_setI2940;
                  end if;
                else
                  \$v2959\ := \$arr1451_ptr_take\;
                  if \$v2959\(0) = '1' then
                    \state\ <= q_wait2958;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
                    \state\ <= pause_setI2956;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811424\;
              end if;
            end if;
          when pause_getII2969 =>
            \$arr1451_ptr_take\(0) := '0';
            \$949_y\ := \$arr1451_value\;
            \$v2966\ := \$arr1452_ptr_take\;
            if \$v2966\(0) = '1' then
              \state\ <= q_wait2965;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2963;
            end if;
          when pause_getII2980 =>
            \$arr1451_ptr_take\(0) := '0';
            \$991\ := \$arr1451_value\;
            \$986\ := \$991\(36 to 71);
            \$v2977\ := \$986\;
            \$v2978\ := \$v2977\(0 to 3);
            \$v2976\ := \$v2977\(4 to 35);
            case \$v2978\ is
            when "0010" =>
              \$987_i\ := \$v2976\(0 to 31);
              \$985\ := \$987_i\;
              if \$984_lock\(0) = '1' then
                \state\ <= get_wait2974;
              else
                \$984_lock\ := eclat_true;
                \state\ <= get_pause2975;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811426\;
            end case;
          when pause_getII2985 =>
            \$arr1452_ptr_take\(0) := '0';
            \$996\ := \$arr1452_value\;
            if \$996_lock\(0) = '1' then
              \state\ <= get_wait2983;
            else
              \$995\ := \$996\;
              \$v2982\ := \$arr1451_ptr_take\;
              if \$v2982\(0) = '1' then
                \state\ <= q_wait2981;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$995\));
                \state\ <= pause_getI2979;
              end if;
            end if;
          when pause_getII2989 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v2987\ := \$arr1452_ptr_take\;
            if \$v2987\(0) = '1' then
              \state\ <= q_wait2986;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2984;
            end if;
          when pause_getII2998 =>
            \$arr1451_ptr_take\(0) := '0';
            \$971\ := \$arr1451_value\;
            \$970\ := \$971\(72 to 107);
            \$v2996\ := "00000000000000000000000000000000";
            \$968\ := "0000" & \$v2996\ & \$969\ & \$970\;
            \$v2995\ := \$arr1451_ptr_take\;
            if \$v2995\(0) = '1' then
              \state\ <= q_wait2994;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$967\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$968\;
              \state\ <= pause_setI2992;
            end if;
          when pause_getII3003 =>
            \$arr1452_ptr_take\(0) := '0';
            \$976\ := \$arr1452_value\;
            if \$976_lock\(0) = '1' then
              \state\ <= get_wait3001;
            else
              \$975\ := \$976\;
              \$v3000\ := \$arr1451_ptr_take\;
              if \$v3000\(0) = '1' then
                \state\ <= q_wait2999;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$975\));
                \state\ <= pause_getI2997;
              end if;
            end if;
          when pause_getII3007 =>
            \$arr1451_ptr_take\(0) := '0';
            \$977\ := \$arr1451_value\;
            \$969\ := \$977\(36 to 71);
            \$v3005\ := \$arr1452_ptr_take\;
            if \$v3005\(0) = '1' then
              \state\ <= q_wait3004;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3002;
            end if;
          when pause_getII3012 =>
            \$arr1452_ptr_take\(0) := '0';
            \$982\ := \$arr1452_value\;
            if \$982_lock\(0) = '1' then
              \state\ <= get_wait3010;
            else
              \$981\ := \$982\;
              \$v3009\ := \$arr1451_ptr_take\;
              if \$v3009\(0) = '1' then
                \state\ <= q_wait3008;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$981\));
                \state\ <= pause_getI3006;
              end if;
            end if;
          when pause_getII3017 =>
            \$arr1452_ptr_take\(0) := '0';
            \$983\ := \$arr1452_value\;
            if \$983_lock\(0) = '1' then
              \state\ <= get_wait3015;
            else
              \$967\ := \$983\;
              \$v3014\ := \$arr1452_ptr_take\;
              if \$v3014\(0) = '1' then
                \state\ <= q_wait3013;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3011;
              end if;
            end if;
          when pause_getII3025 =>
            \$arr1451_ptr_take\(0) := '0';
            \$999\ := \$arr1451_value\;
            \$997\ := \$999\(36 to 71);
            \$v3022\ := \$997\;
            \$v3023\ := \$v3022\(0 to 3);
            \$v3021\ := \$v3022\(4 to 35);
            case \$v3023\ is
            when "0010" =>
              \$966\ := eclat_true;
              \$v3020\ := \$966\;
              if \$v3020\(0) = '1' then
                \$v2991\ := \$arr1452_ptr_take\;
                if \$v2991\(0) = '1' then
                  \state\ <= q_wait2990;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2988;
                end if;
              else
                \$v3019\ := \$arr1452_ptr_take\;
                if \$v3019\(0) = '1' then
                  \state\ <= q_wait3018;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3016;
                end if;
              end if;
            when others =>
              \$966\ := eclat_false;
              \$v3020\ := \$966\;
              if \$v3020\(0) = '1' then
                \$v2991\ := \$arr1452_ptr_take\;
                if \$v2991\(0) = '1' then
                  \state\ <= q_wait2990;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2988;
                end if;
              else
                \$v3019\ := \$arr1452_ptr_take\;
                if \$v3019\(0) = '1' then
                  \state\ <= q_wait3018;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3016;
                end if;
              end if;
            end case;
          when pause_getII3030 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1004\ := \$arr1452_value\;
            if \$1004_lock\(0) = '1' then
              \state\ <= get_wait3028;
            else
              \$1003\ := \$1004\;
              \$v3027\ := \$arr1451_ptr_take\;
              if \$v3027\(0) = '1' then
                \state\ <= q_wait3026;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1003\));
                \state\ <= pause_getI3024;
              end if;
            end if;
          when pause_getII3034 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1005\ := \$arr1451_value\;
            \$965_x\ := \$1005\(0 to 35);
            \$v3032\ := \$arr1452_ptr_take\;
            if \$v3032\(0) = '1' then
              \state\ <= q_wait3031;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3029;
            end if;
          when pause_getII3039 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1010\ := \$arr1452_value\;
            if \$1010_lock\(0) = '1' then
              \state\ <= get_wait3037;
            else
              \$1009\ := \$1010\;
              \$v3036\ := \$arr1451_ptr_take\;
              if \$v3036\(0) = '1' then
                \state\ <= q_wait3035;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1009\));
                \state\ <= pause_getI3033;
              end if;
            end if;
          when pause_getII3048 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1037\ := \$arr1451_value\;
            \$1032\ := \$1037\(36 to 71);
            \$v3045\ := \$1032\;
            \$v3046\ := \$v3045\(0 to 3);
            \$v3044\ := \$v3045\(4 to 35);
            case \$v3046\ is
            when "0010" =>
              \$1033_i\ := \$v3044\(0 to 31);
              \$1031\ := \$1033_i\;
              if \$1030_lock\(0) = '1' then
                \state\ <= get_wait3042;
              else
                \$1030_lock\ := eclat_true;
                \state\ <= get_pause3043;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811427\;
            end case;
          when pause_getII3053 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1042\ := \$arr1452_value\;
            if \$1042_lock\(0) = '1' then
              \state\ <= get_wait3051;
            else
              \$1041\ := \$1042\;
              \$v3050\ := \$arr1451_ptr_take\;
              if \$v3050\(0) = '1' then
                \state\ <= q_wait3049;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1041\));
                \state\ <= pause_getI3047;
              end if;
            end if;
          when pause_getII3057 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3055\ := \$arr1452_ptr_take\;
            if \$v3055\(0) = '1' then
              \state\ <= q_wait3054;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3052;
            end if;
          when pause_getII3066 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1017\ := \$arr1451_value\;
            \$1016\ := \$1017\(72 to 107);
            \$v3064\ := "00000000000000000000000000000000";
            \$1014\ := "0000" & \$v3064\ & \$1015\ & \$1016\;
            \$v3063\ := \$arr1451_ptr_take\;
            if \$v3063\(0) = '1' then
              \state\ <= q_wait3062;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1013\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1014\;
              \state\ <= pause_setI3060;
            end if;
          when pause_getII3071 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1022\ := \$arr1452_value\;
            if \$1022_lock\(0) = '1' then
              \state\ <= get_wait3069;
            else
              \$1021\ := \$1022\;
              \$v3068\ := \$arr1451_ptr_take\;
              if \$v3068\(0) = '1' then
                \state\ <= q_wait3067;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1021\));
                \state\ <= pause_getI3065;
              end if;
            end if;
          when pause_getII3075 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1023\ := \$arr1451_value\;
            \$1015\ := \$1023\(36 to 71);
            \$v3073\ := \$arr1452_ptr_take\;
            if \$v3073\(0) = '1' then
              \state\ <= q_wait3072;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3070;
            end if;
          when pause_getII3080 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1028\ := \$arr1452_value\;
            if \$1028_lock\(0) = '1' then
              \state\ <= get_wait3078;
            else
              \$1027\ := \$1028\;
              \$v3077\ := \$arr1451_ptr_take\;
              if \$v3077\(0) = '1' then
                \state\ <= q_wait3076;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1027\));
                \state\ <= pause_getI3074;
              end if;
            end if;
          when pause_getII3085 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1029\ := \$arr1452_value\;
            if \$1029_lock\(0) = '1' then
              \state\ <= get_wait3083;
            else
              \$1013\ := \$1029\;
              \$v3082\ := \$arr1452_ptr_take\;
              if \$v3082\(0) = '1' then
                \state\ <= q_wait3081;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3079;
              end if;
            end if;
          when pause_getII3093 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1045\ := \$arr1451_value\;
            \$1043\ := \$1045\(36 to 71);
            \$v3090\ := \$1043\;
            \$v3091\ := \$v3090\(0 to 3);
            \$v3089\ := \$v3090\(4 to 35);
            case \$v3091\ is
            when "0010" =>
              \$1012\ := eclat_true;
              \$v3088\ := \$1012\;
              if \$v3088\(0) = '1' then
                \$v3059\ := \$arr1452_ptr_take\;
                if \$v3059\(0) = '1' then
                  \state\ <= q_wait3058;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3056;
                end if;
              else
                \$v3087\ := \$arr1452_ptr_take\;
                if \$v3087\(0) = '1' then
                  \state\ <= q_wait3086;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3084;
                end if;
              end if;
            when others =>
              \$1012\ := eclat_false;
              \$v3088\ := \$1012\;
              if \$v3088\(0) = '1' then
                \$v3059\ := \$arr1452_ptr_take\;
                if \$v3059\(0) = '1' then
                  \state\ <= q_wait3058;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3056;
                end if;
              else
                \$v3087\ := \$arr1452_ptr_take\;
                if \$v3087\(0) = '1' then
                  \state\ <= q_wait3086;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3084;
                end if;
              end if;
            end case;
          when pause_getII3098 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1050\ := \$arr1452_value\;
            if \$1050_lock\(0) = '1' then
              \state\ <= get_wait3096;
            else
              \$1049\ := \$1050\;
              \$v3095\ := \$arr1451_ptr_take\;
              if \$v3095\(0) = '1' then
                \state\ <= q_wait3094;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1049\));
                \state\ <= pause_getI3092;
              end if;
            end if;
          when pause_getII3102 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1051\ := \$arr1451_value\;
            \$1011_x\ := \$1051\(0 to 35);
            \$v3100\ := \$arr1452_ptr_take\;
            if \$v3100\(0) = '1' then
              \state\ <= q_wait3099;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3097;
            end if;
          when pause_getII3107 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1056\ := \$arr1452_value\;
            if \$1056_lock\(0) = '1' then
              \state\ <= get_wait3105;
            else
              \$1055\ := \$1056\;
              \$v3104\ := \$arr1451_ptr_take\;
              if \$v3104\(0) = '1' then
                \state\ <= q_wait3103;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1055\));
                \state\ <= pause_getI3101;
              end if;
            end if;
          when pause_getII3118 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1069\ := \$arr1452_value\;
            if \$1069_lock\(0) = '1' then
              \state\ <= get_wait3116;
            else
              \$1068\ := \$1069\;
              \$1067\ := \$1068\ & "00000000000000000000000000000001";
              \$1066\ := eclat_sub(\$1067\);
              if \$1065_lock\(0) = '1' then
                \state\ <= get_wait3114;
              else
                \$1065_lock\ := eclat_true;
                \state\ <= get_pause3115;
              end if;
            end if;
          when pause_getII3122 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3120\ := \$arr1452_ptr_take\;
            if \$v3120\(0) = '1' then
              \state\ <= q_wait3119;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3117;
            end if;
          when pause_getII3134 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1061_lock\(0) = '1' then
              \state\ <= get_wait3131;
            else
              \$1061_lock\ := eclat_true;
              \state\ <= get_pause3132;
            end if;
          when pause_getII3146 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1073\ := \$arr1452_value\;
            if \$1073_lock\(0) = '1' then
              \state\ <= get_wait3144;
            else
              \$1057_i\ := \$1073\;
              \$v3143\ := eclat_gt(\$1057_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3143\(0) = '1' then
                \$v3142\ := eclat_eq(\$1057_i\ & X"000" & X"15f90");
                if \$v3142\(0) = '1' then
                  \$v3130\ := \$arr1451_ptr_take\;
                  if \$v3130\(0) = '1' then
                    \state\ <= q_wait3129;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3125\ := "00000000000000000000000000000000";
                    \$v3126\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$58_result\(72 to 107) & "0001" & \$v3125\ & "0001" & \$v3126\;
                    \state\ <= pause_setI3127;
                  end if;
                else
                  \$v3141\ := \$arr1451_ptr_take\;
                  if \$v3141\(0) = '1' then
                    \state\ <= q_wait3140;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3137\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$58_result\(72 to 107) & "0010" & \$1057_i\ & "0001" & \$v3137\;
                    \state\ <= pause_setI3138;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811428\;
              end if;
            end if;
          when pause_getII3151 =>
            \$arr1451_ptr_take\(0) := '0';
            \$58_result\ := \$arr1451_value\;
            \$v3148\ := \$arr1452_ptr_take\;
            if \$v3148\(0) = '1' then
              \state\ <= q_wait3147;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3145;
            end if;
          when pause_getII3162 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1105\ := \$arr1451_value\;
            \$1100\ := \$1105\(36 to 71);
            \$v3159\ := \$1100\;
            \$v3160\ := \$v3159\(0 to 3);
            \$v3158\ := \$v3159\(4 to 35);
            case \$v3160\ is
            when "0010" =>
              \$1101_i\ := \$v3158\(0 to 31);
              \$1099\ := \$1101_i\;
              if \$1098_lock\(0) = '1' then
                \state\ <= get_wait3156;
              else
                \$1098_lock\ := eclat_true;
                \state\ <= get_pause3157;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811430\;
            end case;
          when pause_getII3167 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1110\ := \$arr1452_value\;
            if \$1110_lock\(0) = '1' then
              \state\ <= get_wait3165;
            else
              \$1109\ := \$1110\;
              \$v3164\ := \$arr1451_ptr_take\;
              if \$v3164\(0) = '1' then
                \state\ <= q_wait3163;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1109\));
                \state\ <= pause_getI3161;
              end if;
            end if;
          when pause_getII3171 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3169\ := \$arr1452_ptr_take\;
            if \$v3169\(0) = '1' then
              \state\ <= q_wait3168;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3166;
            end if;
          when pause_getII3180 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1085\ := \$arr1451_value\;
            \$1084\ := \$1085\(72 to 107);
            \$v3178\ := "00000000000000000000000000000000";
            \$1082\ := "0000" & \$v3178\ & \$1083\ & \$1084\;
            \$v3177\ := \$arr1451_ptr_take\;
            if \$v3177\(0) = '1' then
              \state\ <= q_wait3176;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1081\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1082\;
              \state\ <= pause_setI3174;
            end if;
          when pause_getII3185 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1090\ := \$arr1452_value\;
            if \$1090_lock\(0) = '1' then
              \state\ <= get_wait3183;
            else
              \$1089\ := \$1090\;
              \$v3182\ := \$arr1451_ptr_take\;
              if \$v3182\(0) = '1' then
                \state\ <= q_wait3181;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1089\));
                \state\ <= pause_getI3179;
              end if;
            end if;
          when pause_getII3189 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1091\ := \$arr1451_value\;
            \$1083\ := \$1091\(36 to 71);
            \$v3187\ := \$arr1452_ptr_take\;
            if \$v3187\(0) = '1' then
              \state\ <= q_wait3186;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3184;
            end if;
          when pause_getII3194 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1096\ := \$arr1452_value\;
            if \$1096_lock\(0) = '1' then
              \state\ <= get_wait3192;
            else
              \$1095\ := \$1096\;
              \$v3191\ := \$arr1451_ptr_take\;
              if \$v3191\(0) = '1' then
                \state\ <= q_wait3190;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1095\));
                \state\ <= pause_getI3188;
              end if;
            end if;
          when pause_getII3199 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1097\ := \$arr1452_value\;
            if \$1097_lock\(0) = '1' then
              \state\ <= get_wait3197;
            else
              \$1081\ := \$1097\;
              \$v3196\ := \$arr1452_ptr_take\;
              if \$v3196\(0) = '1' then
                \state\ <= q_wait3195;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3193;
              end if;
            end if;
          when pause_getII3207 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1113\ := \$arr1451_value\;
            \$1111\ := \$1113\(36 to 71);
            \$v3204\ := \$1111\;
            \$v3205\ := \$v3204\(0 to 3);
            \$v3203\ := \$v3204\(4 to 35);
            case \$v3205\ is
            when "0010" =>
              \$1080\ := eclat_true;
              \$v3202\ := \$1080\;
              if \$v3202\(0) = '1' then
                \$v3173\ := \$arr1452_ptr_take\;
                if \$v3173\(0) = '1' then
                  \state\ <= q_wait3172;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3170;
                end if;
              else
                \$v3201\ := \$arr1452_ptr_take\;
                if \$v3201\(0) = '1' then
                  \state\ <= q_wait3200;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3198;
                end if;
              end if;
            when others =>
              \$1080\ := eclat_false;
              \$v3202\ := \$1080\;
              if \$v3202\(0) = '1' then
                \$v3173\ := \$arr1452_ptr_take\;
                if \$v3173\(0) = '1' then
                  \state\ <= q_wait3172;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3170;
                end if;
              else
                \$v3201\ := \$arr1452_ptr_take\;
                if \$v3201\(0) = '1' then
                  \state\ <= q_wait3200;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3198;
                end if;
              end if;
            end case;
          when pause_getII3212 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1118\ := \$arr1452_value\;
            if \$1118_lock\(0) = '1' then
              \state\ <= get_wait3210;
            else
              \$1117\ := \$1118\;
              \$v3209\ := \$arr1451_ptr_take\;
              if \$v3209\(0) = '1' then
                \state\ <= q_wait3208;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1117\));
                \state\ <= pause_getI3206;
              end if;
            end if;
          when pause_getII3216 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1119\ := \$arr1451_value\;
            \$1079_x\ := \$1119\(0 to 35);
            \$v3214\ := \$arr1452_ptr_take\;
            if \$v3214\(0) = '1' then
              \state\ <= q_wait3213;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3211;
            end if;
          when pause_getII3221 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1124\ := \$arr1452_value\;
            if \$1124_lock\(0) = '1' then
              \state\ <= get_wait3219;
            else
              \$1123\ := \$1124\;
              \$v3218\ := \$arr1451_ptr_take\;
              if \$v3218\(0) = '1' then
                \state\ <= q_wait3217;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1123\));
                \state\ <= pause_getI3215;
              end if;
            end if;
          when pause_getII3232 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1138\ := \$arr1452_value\;
            if \$1138_lock\(0) = '1' then
              \state\ <= get_wait3230;
            else
              \$1137\ := \$1138\;
              \$1136\ := \$1137\ & "00000000000000000000000000000001";
              \$1135\ := eclat_sub(\$1136\);
              if \$1134_lock\(0) = '1' then
                \state\ <= get_wait3228;
              else
                \$1134_lock\ := eclat_true;
                \state\ <= get_pause3229;
              end if;
            end if;
          when pause_getII3236 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3234\ := \$arr1452_ptr_take\;
            if \$v3234\(0) = '1' then
              \state\ <= q_wait3233;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3231;
            end if;
          when pause_getII3248 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1130_lock\(0) = '1' then
              \state\ <= get_wait3245;
            else
              \$1130_lock\ := eclat_true;
              \state\ <= get_pause3246;
            end if;
          when pause_getII3260 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1142\ := \$arr1452_value\;
            if \$1142_lock\(0) = '1' then
              \state\ <= get_wait3258;
            else
              \$1126_i\ := \$1142\;
              \$v3257\ := eclat_gt(\$1126_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3257\(0) = '1' then
                \$v3256\ := eclat_eq(\$1126_i\ & X"000" & X"15f90");
                if \$v3256\(0) = '1' then
                  \$v3244\ := \$arr1451_ptr_take\;
                  if \$v3244\(0) = '1' then
                    \state\ <= q_wait3243;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3239\ := "00000000000000000000000000000000";
                    \$v3240\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1125_result\(36 to 71) & "0001" & \$v3239\ & "0001" & \$v3240\;
                    \state\ <= pause_setI3241;
                  end if;
                else
                  \$v3255\ := \$arr1451_ptr_take\;
                  if \$v3255\(0) = '1' then
                    \state\ <= q_wait3254;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3251\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1125_result\(36 to 71) & "0010" & \$1126_i\ & "0001" & \$v3251\;
                    \state\ <= pause_setI3252;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811431\;
              end if;
            end if;
          when pause_getII3265 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1125_result\ := \$arr1451_value\;
            \$v3262\ := \$arr1452_ptr_take\;
            if \$v3262\(0) = '1' then
              \state\ <= q_wait3261;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3259;
            end if;
          when pause_getII3276 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1174\ := \$arr1451_value\;
            \$1169\ := \$1174\(36 to 71);
            \$v3273\ := \$1169\;
            \$v3274\ := \$v3273\(0 to 3);
            \$v3272\ := \$v3273\(4 to 35);
            case \$v3274\ is
            when "0010" =>
              \$1170_i\ := \$v3272\(0 to 31);
              \$1168\ := \$1170_i\;
              if \$1167_lock\(0) = '1' then
                \state\ <= get_wait3270;
              else
                \$1167_lock\ := eclat_true;
                \state\ <= get_pause3271;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811433\;
            end case;
          when pause_getII3281 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1179\ := \$arr1452_value\;
            if \$1179_lock\(0) = '1' then
              \state\ <= get_wait3279;
            else
              \$1178\ := \$1179\;
              \$v3278\ := \$arr1451_ptr_take\;
              if \$v3278\(0) = '1' then
                \state\ <= q_wait3277;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1178\));
                \state\ <= pause_getI3275;
              end if;
            end if;
          when pause_getII3285 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3283\ := \$arr1452_ptr_take\;
            if \$v3283\(0) = '1' then
              \state\ <= q_wait3282;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3280;
            end if;
          when pause_getII3294 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1154\ := \$arr1451_value\;
            \$1153\ := \$1154\(72 to 107);
            \$v3292\ := "00000000000000000000000000000000";
            \$1151\ := "0000" & \$v3292\ & \$1152\ & \$1153\;
            \$v3291\ := \$arr1451_ptr_take\;
            if \$v3291\(0) = '1' then
              \state\ <= q_wait3290;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1150\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1151\;
              \state\ <= pause_setI3288;
            end if;
          when pause_getII3299 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1159\ := \$arr1452_value\;
            if \$1159_lock\(0) = '1' then
              \state\ <= get_wait3297;
            else
              \$1158\ := \$1159\;
              \$v3296\ := \$arr1451_ptr_take\;
              if \$v3296\(0) = '1' then
                \state\ <= q_wait3295;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1158\));
                \state\ <= pause_getI3293;
              end if;
            end if;
          when pause_getII3303 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1160\ := \$arr1451_value\;
            \$1152\ := \$1160\(36 to 71);
            \$v3301\ := \$arr1452_ptr_take\;
            if \$v3301\(0) = '1' then
              \state\ <= q_wait3300;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3298;
            end if;
          when pause_getII3308 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1165\ := \$arr1452_value\;
            if \$1165_lock\(0) = '1' then
              \state\ <= get_wait3306;
            else
              \$1164\ := \$1165\;
              \$v3305\ := \$arr1451_ptr_take\;
              if \$v3305\(0) = '1' then
                \state\ <= q_wait3304;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1164\));
                \state\ <= pause_getI3302;
              end if;
            end if;
          when pause_getII3313 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1166\ := \$arr1452_value\;
            if \$1166_lock\(0) = '1' then
              \state\ <= get_wait3311;
            else
              \$1150\ := \$1166\;
              \$v3310\ := \$arr1452_ptr_take\;
              if \$v3310\(0) = '1' then
                \state\ <= q_wait3309;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3307;
              end if;
            end if;
          when pause_getII3321 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1182\ := \$arr1451_value\;
            \$1180\ := \$1182\(36 to 71);
            \$v3318\ := \$1180\;
            \$v3319\ := \$v3318\(0 to 3);
            \$v3317\ := \$v3318\(4 to 35);
            case \$v3319\ is
            when "0010" =>
              \$1149\ := eclat_true;
              \$v3316\ := \$1149\;
              if \$v3316\(0) = '1' then
                \$v3287\ := \$arr1452_ptr_take\;
                if \$v3287\(0) = '1' then
                  \state\ <= q_wait3286;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3284;
                end if;
              else
                \$v3315\ := \$arr1452_ptr_take\;
                if \$v3315\(0) = '1' then
                  \state\ <= q_wait3314;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3312;
                end if;
              end if;
            when others =>
              \$1149\ := eclat_false;
              \$v3316\ := \$1149\;
              if \$v3316\(0) = '1' then
                \$v3287\ := \$arr1452_ptr_take\;
                if \$v3287\(0) = '1' then
                  \state\ <= q_wait3286;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3284;
                end if;
              else
                \$v3315\ := \$arr1452_ptr_take\;
                if \$v3315\(0) = '1' then
                  \state\ <= q_wait3314;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3312;
                end if;
              end if;
            end case;
          when pause_getII3326 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1187\ := \$arr1452_value\;
            if \$1187_lock\(0) = '1' then
              \state\ <= get_wait3324;
            else
              \$1186\ := \$1187\;
              \$v3323\ := \$arr1451_ptr_take\;
              if \$v3323\(0) = '1' then
                \state\ <= q_wait3322;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1186\));
                \state\ <= pause_getI3320;
              end if;
            end if;
          when pause_getII3330 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1188\ := \$arr1451_value\;
            \$1148_x\ := \$1188\(0 to 35);
            \$v3328\ := \$arr1452_ptr_take\;
            if \$v3328\(0) = '1' then
              \state\ <= q_wait3327;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3325;
            end if;
          when pause_getII3335 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1193\ := \$arr1452_value\;
            if \$1193_lock\(0) = '1' then
              \state\ <= get_wait3333;
            else
              \$1192\ := \$1193\;
              \$v3332\ := \$arr1451_ptr_take\;
              if \$v3332\(0) = '1' then
                \state\ <= q_wait3331;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1192\));
                \state\ <= pause_getI3329;
              end if;
            end if;
          when pause_getII3346 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1207\ := \$arr1452_value\;
            if \$1207_lock\(0) = '1' then
              \state\ <= get_wait3344;
            else
              \$1206\ := \$1207\;
              \$1205\ := \$1206\ & "00000000000000000000000000000001";
              \$1204\ := eclat_sub(\$1205\);
              if \$1203_lock\(0) = '1' then
                \state\ <= get_wait3342;
              else
                \$1203_lock\ := eclat_true;
                \state\ <= get_pause3343;
              end if;
            end if;
          when pause_getII3350 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3348\ := \$arr1452_ptr_take\;
            if \$v3348\(0) = '1' then
              \state\ <= q_wait3347;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3345;
            end if;
          when pause_getII3362 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1199_lock\(0) = '1' then
              \state\ <= get_wait3359;
            else
              \$1199_lock\ := eclat_true;
              \state\ <= get_pause3360;
            end if;
          when pause_getII3374 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1211\ := \$arr1452_value\;
            if \$1211_lock\(0) = '1' then
              \state\ <= get_wait3372;
            else
              \$1195_i\ := \$1211\;
              \$v3371\ := eclat_gt(\$1195_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3371\(0) = '1' then
                \$v3370\ := eclat_eq(\$1195_i\ & X"000" & X"15f90");
                if \$v3370\(0) = '1' then
                  \$v3358\ := \$arr1451_ptr_take\;
                  if \$v3358\(0) = '1' then
                    \state\ <= q_wait3357;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3353\ := "00000000000000000000000000000000";
                    \$v3354\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1194_result\(0 to 35) & "0001" & \$v3353\ & "0001" & \$v3354\;
                    \state\ <= pause_setI3355;
                  end if;
                else
                  \$v3369\ := \$arr1451_ptr_take\;
                  if \$v3369\(0) = '1' then
                    \state\ <= q_wait3368;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3365\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1194_result\(0 to 35) & "0010" & \$1195_i\ & "0001" & \$v3365\;
                    \state\ <= pause_setI3366;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811434\;
              end if;
            end if;
          when pause_getII3379 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1194_result\ := \$arr1451_value\;
            \$v3376\ := \$arr1452_ptr_take\;
            if \$v3376\(0) = '1' then
              \state\ <= q_wait3375;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3373;
            end if;
          when pause_getII3390 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1243\ := \$arr1451_value\;
            \$1238\ := \$1243\(36 to 71);
            \$v3387\ := \$1238\;
            \$v3388\ := \$v3387\(0 to 3);
            \$v3386\ := \$v3387\(4 to 35);
            case \$v3388\ is
            when "0010" =>
              \$1239_i\ := \$v3386\(0 to 31);
              \$1237\ := \$1239_i\;
              if \$1236_lock\(0) = '1' then
                \state\ <= get_wait3384;
              else
                \$1236_lock\ := eclat_true;
                \state\ <= get_pause3385;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811436\;
            end case;
          when pause_getII3395 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1248\ := \$arr1452_value\;
            if \$1248_lock\(0) = '1' then
              \state\ <= get_wait3393;
            else
              \$1247\ := \$1248\;
              \$v3392\ := \$arr1451_ptr_take\;
              if \$v3392\(0) = '1' then
                \state\ <= q_wait3391;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1247\));
                \state\ <= pause_getI3389;
              end if;
            end if;
          when pause_getII3399 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3397\ := \$arr1452_ptr_take\;
            if \$v3397\(0) = '1' then
              \state\ <= q_wait3396;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3394;
            end if;
          when pause_getII3408 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1223\ := \$arr1451_value\;
            \$1222\ := \$1223\(72 to 107);
            \$v3406\ := "00000000000000000000000000000000";
            \$1220\ := "0000" & \$v3406\ & \$1221\ & \$1222\;
            \$v3405\ := \$arr1451_ptr_take\;
            if \$v3405\(0) = '1' then
              \state\ <= q_wait3404;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1219\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1220\;
              \state\ <= pause_setI3402;
            end if;
          when pause_getII3413 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1228\ := \$arr1452_value\;
            if \$1228_lock\(0) = '1' then
              \state\ <= get_wait3411;
            else
              \$1227\ := \$1228\;
              \$v3410\ := \$arr1451_ptr_take\;
              if \$v3410\(0) = '1' then
                \state\ <= q_wait3409;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1227\));
                \state\ <= pause_getI3407;
              end if;
            end if;
          when pause_getII3417 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1229\ := \$arr1451_value\;
            \$1221\ := \$1229\(36 to 71);
            \$v3415\ := \$arr1452_ptr_take\;
            if \$v3415\(0) = '1' then
              \state\ <= q_wait3414;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3412;
            end if;
          when pause_getII3422 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1234\ := \$arr1452_value\;
            if \$1234_lock\(0) = '1' then
              \state\ <= get_wait3420;
            else
              \$1233\ := \$1234\;
              \$v3419\ := \$arr1451_ptr_take\;
              if \$v3419\(0) = '1' then
                \state\ <= q_wait3418;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1233\));
                \state\ <= pause_getI3416;
              end if;
            end if;
          when pause_getII3427 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1235\ := \$arr1452_value\;
            if \$1235_lock\(0) = '1' then
              \state\ <= get_wait3425;
            else
              \$1219\ := \$1235\;
              \$v3424\ := \$arr1452_ptr_take\;
              if \$v3424\(0) = '1' then
                \state\ <= q_wait3423;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3421;
              end if;
            end if;
          when pause_getII3435 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1251\ := \$arr1451_value\;
            \$1249\ := \$1251\(36 to 71);
            \$v3432\ := \$1249\;
            \$v3433\ := \$v3432\(0 to 3);
            \$v3431\ := \$v3432\(4 to 35);
            case \$v3433\ is
            when "0010" =>
              \$1218\ := eclat_true;
              \$v3430\ := \$1218\;
              if \$v3430\(0) = '1' then
                \$v3401\ := \$arr1452_ptr_take\;
                if \$v3401\(0) = '1' then
                  \state\ <= q_wait3400;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3398;
                end if;
              else
                \$v3429\ := \$arr1452_ptr_take\;
                if \$v3429\(0) = '1' then
                  \state\ <= q_wait3428;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3426;
                end if;
              end if;
            when others =>
              \$1218\ := eclat_false;
              \$v3430\ := \$1218\;
              if \$v3430\(0) = '1' then
                \$v3401\ := \$arr1452_ptr_take\;
                if \$v3401\(0) = '1' then
                  \state\ <= q_wait3400;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3398;
                end if;
              else
                \$v3429\ := \$arr1452_ptr_take\;
                if \$v3429\(0) = '1' then
                  \state\ <= q_wait3428;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3426;
                end if;
              end if;
            end case;
          when pause_getII3440 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1256\ := \$arr1452_value\;
            if \$1256_lock\(0) = '1' then
              \state\ <= get_wait3438;
            else
              \$1255\ := \$1256\;
              \$v3437\ := \$arr1451_ptr_take\;
              if \$v3437\(0) = '1' then
                \state\ <= q_wait3436;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1255\));
                \state\ <= pause_getI3434;
              end if;
            end if;
          when pause_getII3444 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1257\ := \$arr1451_value\;
            \$1217_x\ := \$1257\(0 to 35);
            \$v3442\ := \$arr1452_ptr_take\;
            if \$v3442\(0) = '1' then
              \state\ <= q_wait3441;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3439;
            end if;
          when pause_getII3449 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1262\ := \$arr1452_value\;
            if \$1262_lock\(0) = '1' then
              \state\ <= get_wait3447;
            else
              \$1261\ := \$1262\;
              \$v3446\ := \$arr1451_ptr_take\;
              if \$v3446\(0) = '1' then
                \state\ <= q_wait3445;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1261\));
                \state\ <= pause_getI3443;
              end if;
            end if;
          when pause_getII3459 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1268_lock\(0) = '1' then
              \state\ <= get_wait3456;
            else
              \$1268_lock\ := eclat_true;
              \state\ <= get_pause3457;
            end if;
          when pause_getII3469 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1267_lock\(0) = '1' then
              \state\ <= get_wait3466;
            else
              \$1267_lock\ := eclat_true;
              \state\ <= get_pause3467;
            end if;
          when pause_getII3486 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1269\ := \$arr1452_value\;
            if \$1269_lock\(0) = '1' then
              \state\ <= get_wait3484;
            else
              \$1263_i\ := \$1269\;
              \$v3483\ := eclat_gt(\$1263_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3483\(0) = '1' then
                \$v3482\ := eclat_eq(\$1263_i\ & X"000" & X"15f90");
                if \$v3482\(0) = '1' then
                  \$v3465\ := \$arr1451_ptr_take\;
                  if \$v3465\(0) = '1' then
                    \state\ <= q_wait3464;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$74_result_after_f\;
                    \state\ <= pause_setI3462;
                  end if;
                else
                  \$v3481\ := \$arr1451_ptr_take\;
                  if \$v3481\(0) = '1' then
                    \state\ <= q_wait3480;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$74_result_after_f\;
                    \state\ <= pause_setI3478;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811437\;
              end if;
            end if;
          when pause_getII3504 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1296\ := \$arr1451_value\;
            \$1291\ := \$1296\(36 to 71);
            \$v3501\ := \$1291\;
            \$v3502\ := \$v3501\(0 to 3);
            \$v3500\ := \$v3501\(4 to 35);
            case \$v3502\ is
            when "0010" =>
              \$1292_i\ := \$v3500\(0 to 31);
              \$1290\ := \$1292_i\;
              if \$1289_lock\(0) = '1' then
                \state\ <= get_wait3498;
              else
                \$1289_lock\ := eclat_true;
                \state\ <= get_pause3499;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811438\;
            end case;
          when pause_getII3509 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1301\ := \$arr1452_value\;
            if \$1301_lock\(0) = '1' then
              \state\ <= get_wait3507;
            else
              \$1300\ := \$1301\;
              \$v3506\ := \$arr1451_ptr_take\;
              if \$v3506\(0) = '1' then
                \state\ <= q_wait3505;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1300\));
                \state\ <= pause_getI3503;
              end if;
            end if;
          when pause_getII3513 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3511\ := \$arr1452_ptr_take\;
            if \$v3511\(0) = '1' then
              \state\ <= q_wait3510;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3508;
            end if;
          when pause_getII3522 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1276\ := \$arr1451_value\;
            \$1275\ := \$1276\(72 to 107);
            \$v3520\ := "00000000000000000000000000000000";
            \$1273\ := "0000" & \$v3520\ & \$1274\ & \$1275\;
            \$v3519\ := \$arr1451_ptr_take\;
            if \$v3519\(0) = '1' then
              \state\ <= q_wait3518;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1272\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1273\;
              \state\ <= pause_setI3516;
            end if;
          when pause_getII3527 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1281\ := \$arr1452_value\;
            if \$1281_lock\(0) = '1' then
              \state\ <= get_wait3525;
            else
              \$1280\ := \$1281\;
              \$v3524\ := \$arr1451_ptr_take\;
              if \$v3524\(0) = '1' then
                \state\ <= q_wait3523;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1280\));
                \state\ <= pause_getI3521;
              end if;
            end if;
          when pause_getII3531 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1282\ := \$arr1451_value\;
            \$1274\ := \$1282\(36 to 71);
            \$v3529\ := \$arr1452_ptr_take\;
            if \$v3529\(0) = '1' then
              \state\ <= q_wait3528;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3526;
            end if;
          when pause_getII3536 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1287\ := \$arr1452_value\;
            if \$1287_lock\(0) = '1' then
              \state\ <= get_wait3534;
            else
              \$1286\ := \$1287\;
              \$v3533\ := \$arr1451_ptr_take\;
              if \$v3533\(0) = '1' then
                \state\ <= q_wait3532;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1286\));
                \state\ <= pause_getI3530;
              end if;
            end if;
          when pause_getII3541 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1288\ := \$arr1452_value\;
            if \$1288_lock\(0) = '1' then
              \state\ <= get_wait3539;
            else
              \$1272\ := \$1288\;
              \$v3538\ := \$arr1452_ptr_take\;
              if \$v3538\(0) = '1' then
                \state\ <= q_wait3537;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3535;
              end if;
            end if;
          when pause_getII3549 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1304\ := \$arr1451_value\;
            \$1302\ := \$1304\(36 to 71);
            \$v3546\ := \$1302\;
            \$v3547\ := \$v3546\(0 to 3);
            \$v3545\ := \$v3546\(4 to 35);
            case \$v3547\ is
            when "0010" =>
              \$1271\ := eclat_true;
              \$v3544\ := \$1271\;
              if \$v3544\(0) = '1' then
                \$v3515\ := \$arr1452_ptr_take\;
                if \$v3515\(0) = '1' then
                  \state\ <= q_wait3514;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3512;
                end if;
              else
                \$v3543\ := \$arr1452_ptr_take\;
                if \$v3543\(0) = '1' then
                  \state\ <= q_wait3542;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3540;
                end if;
              end if;
            when others =>
              \$1271\ := eclat_false;
              \$v3544\ := \$1271\;
              if \$v3544\(0) = '1' then
                \$v3515\ := \$arr1452_ptr_take\;
                if \$v3515\(0) = '1' then
                  \state\ <= q_wait3514;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3512;
                end if;
              else
                \$v3543\ := \$arr1452_ptr_take\;
                if \$v3543\(0) = '1' then
                  \state\ <= q_wait3542;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3540;
                end if;
              end if;
            end case;
          when pause_getII3554 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1309\ := \$arr1452_value\;
            if \$1309_lock\(0) = '1' then
              \state\ <= get_wait3552;
            else
              \$1308\ := \$1309\;
              \$v3551\ := \$arr1451_ptr_take\;
              if \$v3551\(0) = '1' then
                \state\ <= q_wait3550;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1308\));
                \state\ <= pause_getI3548;
              end if;
            end if;
          when pause_getII3558 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1310\ := \$arr1451_value\;
            \$1270_x\ := \$1310\(0 to 35);
            \$v3556\ := \$arr1452_ptr_take\;
            if \$v3556\(0) = '1' then
              \state\ <= q_wait3555;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3553;
            end if;
          when pause_getII3563 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1315\ := \$arr1452_value\;
            if \$1315_lock\(0) = '1' then
              \state\ <= get_wait3561;
            else
              \$1314\ := \$1315\;
              \$v3560\ := \$arr1451_ptr_take\;
              if \$v3560\(0) = '1' then
                \state\ <= q_wait3559;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1314\));
                \state\ <= pause_getI3557;
              end if;
            end if;
          when pause_getII3573 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1324_lock\(0) = '1' then
              \state\ <= get_wait3570;
            else
              \$1324_lock\ := eclat_true;
              \state\ <= get_pause3571;
            end if;
          when pause_getII3584 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1320_lock\(0) = '1' then
              \state\ <= get_wait3581;
            else
              \$1320_lock\ := eclat_true;
              \state\ <= get_pause3582;
            end if;
          when pause_getII3602 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1328\ := \$arr1452_value\;
            if \$1328_lock\(0) = '1' then
              \state\ <= get_wait3600;
            else
              \$1316_i\ := \$1328\;
              \$v3599\ := eclat_gt(\$1316_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3599\(0) = '1' then
                \$v3598\ := eclat_eq(\$1316_i\ & X"000" & X"15f90");
                if \$v3598\(0) = '1' then
                  \$v3580\ := \$arr1451_ptr_take\;
                  if \$v3580\(0) = '1' then
                    \state\ <= q_wait3579;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3576\ := "00000000000000000000000000000001";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3576\;
                    \state\ <= pause_setI3577;
                  end if;
                else
                  \$v3597\ := \$arr1451_ptr_take\;
                  if \$v3597\(0) = '1' then
                    \state\ <= q_wait3596;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3593\ := "00000000000000000000000000000001";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3593\;
                    \state\ <= pause_setI3594;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811439\;
              end if;
            end if;
          when pause_getII3606 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v80\ := \$arr1451_value\;
            \$61_y\ := \$v80\(36 to 71);
            \$v3604\ := \$arr1452_ptr_take\;
            if \$v3604\(0) = '1' then
              \state\ <= q_wait3603;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3601;
            end if;
          when pause_getII3611 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v78\ := \$arr1452_value\;
            if \$v78_lock\(0) = '1' then
              \state\ <= get_wait3609;
            else
              \$v79\ := \$v78\;
              \$v3608\ := \$arr1451_ptr_take\;
              if \$v3608\(0) = '1' then
                \state\ <= q_wait3607;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v79\));
                \state\ <= pause_getI3605;
              end if;
            end if;
          when pause_getII3616 =>
            \$arr1451_ptr_take\(0) := '0';
            \$59_tos\ := \$arr1451_value\;
            \$v3613\ := \$arr1452_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3610;
            end if;
          when pause_getII3627 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1363\ := \$arr1451_value\;
            \$1358\ := \$1363\(36 to 71);
            \$v3624\ := \$1358\;
            \$v3625\ := \$v3624\(0 to 3);
            \$v3623\ := \$v3624\(4 to 35);
            case \$v3625\ is
            when "0010" =>
              \$1359_i\ := \$v3623\(0 to 31);
              \$1357\ := \$1359_i\;
              if \$1356_lock\(0) = '1' then
                \state\ <= get_wait3621;
              else
                \$1356_lock\ := eclat_true;
                \state\ <= get_pause3622;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811441\;
            end case;
          when pause_getII3632 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1368\ := \$arr1452_value\;
            if \$1368_lock\(0) = '1' then
              \state\ <= get_wait3630;
            else
              \$1367\ := \$1368\;
              \$v3629\ := \$arr1451_ptr_take\;
              if \$v3629\(0) = '1' then
                \state\ <= q_wait3628;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1367\));
                \state\ <= pause_getI3626;
              end if;
            end if;
          when pause_getII3636 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3634\ := \$arr1452_ptr_take\;
            if \$v3634\(0) = '1' then
              \state\ <= q_wait3633;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3631;
            end if;
          when pause_getII3645 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1343\ := \$arr1451_value\;
            \$1342\ := \$1343\(72 to 107);
            \$v3643\ := "00000000000000000000000000000000";
            \$1340\ := "0000" & \$v3643\ & \$1341\ & \$1342\;
            \$v3642\ := \$arr1451_ptr_take\;
            if \$v3642\(0) = '1' then
              \state\ <= q_wait3641;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1339\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1340\;
              \state\ <= pause_setI3639;
            end if;
          when pause_getII3650 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1348\ := \$arr1452_value\;
            if \$1348_lock\(0) = '1' then
              \state\ <= get_wait3648;
            else
              \$1347\ := \$1348\;
              \$v3647\ := \$arr1451_ptr_take\;
              if \$v3647\(0) = '1' then
                \state\ <= q_wait3646;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1347\));
                \state\ <= pause_getI3644;
              end if;
            end if;
          when pause_getII3654 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1349\ := \$arr1451_value\;
            \$1341\ := \$1349\(36 to 71);
            \$v3652\ := \$arr1452_ptr_take\;
            if \$v3652\(0) = '1' then
              \state\ <= q_wait3651;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3649;
            end if;
          when pause_getII3659 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1354\ := \$arr1452_value\;
            if \$1354_lock\(0) = '1' then
              \state\ <= get_wait3657;
            else
              \$1353\ := \$1354\;
              \$v3656\ := \$arr1451_ptr_take\;
              if \$v3656\(0) = '1' then
                \state\ <= q_wait3655;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1353\));
                \state\ <= pause_getI3653;
              end if;
            end if;
          when pause_getII3664 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1355\ := \$arr1452_value\;
            if \$1355_lock\(0) = '1' then
              \state\ <= get_wait3662;
            else
              \$1339\ := \$1355\;
              \$v3661\ := \$arr1452_ptr_take\;
              if \$v3661\(0) = '1' then
                \state\ <= q_wait3660;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3658;
              end if;
            end if;
          when pause_getII3672 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1371\ := \$arr1451_value\;
            \$1369\ := \$1371\(36 to 71);
            \$v3669\ := \$1369\;
            \$v3670\ := \$v3669\(0 to 3);
            \$v3668\ := \$v3669\(4 to 35);
            case \$v3670\ is
            when "0010" =>
              \$1338\ := eclat_true;
              \$v3667\ := \$1338\;
              if \$v3667\(0) = '1' then
                \$v3638\ := \$arr1452_ptr_take\;
                if \$v3638\(0) = '1' then
                  \state\ <= q_wait3637;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3635;
                end if;
              else
                \$v3666\ := \$arr1452_ptr_take\;
                if \$v3666\(0) = '1' then
                  \state\ <= q_wait3665;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3663;
                end if;
              end if;
            when others =>
              \$1338\ := eclat_false;
              \$v3667\ := \$1338\;
              if \$v3667\(0) = '1' then
                \$v3638\ := \$arr1452_ptr_take\;
                if \$v3638\(0) = '1' then
                  \state\ <= q_wait3637;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3635;
                end if;
              else
                \$v3666\ := \$arr1452_ptr_take\;
                if \$v3666\(0) = '1' then
                  \state\ <= q_wait3665;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3663;
                end if;
              end if;
            end case;
          when pause_getII3677 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1376\ := \$arr1452_value\;
            if \$1376_lock\(0) = '1' then
              \state\ <= get_wait3675;
            else
              \$1375\ := \$1376\;
              \$v3674\ := \$arr1451_ptr_take\;
              if \$v3674\(0) = '1' then
                \state\ <= q_wait3673;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1375\));
                \state\ <= pause_getI3671;
              end if;
            end if;
          when pause_getII3681 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1377\ := \$arr1451_value\;
            \$1337_x\ := \$1377\(0 to 35);
            \$v3679\ := \$arr1452_ptr_take\;
            if \$v3679\(0) = '1' then
              \state\ <= q_wait3678;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3676;
            end if;
          when pause_getII3686 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1382\ := \$arr1452_value\;
            if \$1382_lock\(0) = '1' then
              \state\ <= get_wait3684;
            else
              \$1381\ := \$1382\;
              \$v3683\ := \$arr1451_ptr_take\;
              if \$v3683\(0) = '1' then
                \state\ <= q_wait3682;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1381\));
                \state\ <= pause_getI3680;
              end if;
            end if;
          when pause_getII3697 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1394\ := \$arr1452_value\;
            if \$1394_lock\(0) = '1' then
              \state\ <= get_wait3695;
            else
              \$1393\ := \$1394\;
              \$1392\ := \$1393\ & "00000000000000000000000000000001";
              \$1391\ := eclat_sub(\$1392\);
              if \$1390_lock\(0) = '1' then
                \state\ <= get_wait3693;
              else
                \$1390_lock\ := eclat_true;
                \state\ <= get_pause3694;
              end if;
            end if;
          when pause_getII3701 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3699\ := \$arr1452_ptr_take\;
            if \$v3699\(0) = '1' then
              \state\ <= q_wait3698;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3696;
            end if;
          when pause_getII3713 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1389_lock\(0) = '1' then
              \state\ <= get_wait3710;
            else
              \$1389_lock\ := eclat_true;
              \state\ <= get_pause3711;
            end if;
          when pause_getII3725 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1395\ := \$arr1452_value\;
            if \$1395_lock\(0) = '1' then
              \state\ <= get_wait3723;
            else
              \$1385_i\ := \$1395\;
              \$v3722\ := eclat_gt(\$1385_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3722\(0) = '1' then
                \$v3721\ := eclat_eq(\$1385_i\ & X"000" & X"15f90");
                if \$v3721\(0) = '1' then
                  \$v3709\ := \$arr1451_ptr_take\;
                  if \$v3709\(0) = '1' then
                    \state\ <= q_wait3708;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3704\ := "00000000000000000000000000000000";
                    \$v3705\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1383_x\ & "0001" & \$v3704\ & "0001" & \$v3705\;
                    \state\ <= pause_setI3706;
                  end if;
                else
                  \$v3720\ := \$arr1451_ptr_take\;
                  if \$v3720\(0) = '1' then
                    \state\ <= q_wait3719;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3716\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$1383_x\ & "0010" & \$1385_i\ & "0001" & \$v3716\;
                    \state\ <= pause_setI3717;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811442\;
              end if;
            end if;
          when pause_getII3734 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1422\ := \$arr1451_value\;
            \$1417\ := \$1422\(36 to 71);
            \$v3731\ := \$1417\;
            \$v3732\ := \$v3731\(0 to 3);
            \$v3730\ := \$v3731\(4 to 35);
            case \$v3732\ is
            when "0010" =>
              \$1418_i\ := \$v3730\(0 to 31);
              \$1416\ := \$1418_i\;
              if \$1415_lock\(0) = '1' then
                \state\ <= get_wait3728;
              else
                \$1415_lock\ := eclat_true;
                \state\ <= get_pause3729;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811443\;
            end case;
          when pause_getII3739 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1427\ := \$arr1452_value\;
            if \$1427_lock\(0) = '1' then
              \state\ <= get_wait3737;
            else
              \$1426\ := \$1427\;
              \$v3736\ := \$arr1451_ptr_take\;
              if \$v3736\(0) = '1' then
                \state\ <= q_wait3735;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1426\));
                \state\ <= pause_getI3733;
              end if;
            end if;
          when pause_getII3743 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3741\ := \$arr1452_ptr_take\;
            if \$v3741\(0) = '1' then
              \state\ <= q_wait3740;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3738;
            end if;
          when pause_getII3752 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1402\ := \$arr1451_value\;
            \$1401\ := \$1402\(72 to 107);
            \$v3750\ := "00000000000000000000000000000000";
            \$1399\ := "0000" & \$v3750\ & \$1400\ & \$1401\;
            \$v3749\ := \$arr1451_ptr_take\;
            if \$v3749\(0) = '1' then
              \state\ <= q_wait3748;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1398\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1399\;
              \state\ <= pause_setI3746;
            end if;
          when pause_getII3757 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1407\ := \$arr1452_value\;
            if \$1407_lock\(0) = '1' then
              \state\ <= get_wait3755;
            else
              \$1406\ := \$1407\;
              \$v3754\ := \$arr1451_ptr_take\;
              if \$v3754\(0) = '1' then
                \state\ <= q_wait3753;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1406\));
                \state\ <= pause_getI3751;
              end if;
            end if;
          when pause_getII3761 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1408\ := \$arr1451_value\;
            \$1400\ := \$1408\(36 to 71);
            \$v3759\ := \$arr1452_ptr_take\;
            if \$v3759\(0) = '1' then
              \state\ <= q_wait3758;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3756;
            end if;
          when pause_getII3766 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1413\ := \$arr1452_value\;
            if \$1413_lock\(0) = '1' then
              \state\ <= get_wait3764;
            else
              \$1412\ := \$1413\;
              \$v3763\ := \$arr1451_ptr_take\;
              if \$v3763\(0) = '1' then
                \state\ <= q_wait3762;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1412\));
                \state\ <= pause_getI3760;
              end if;
            end if;
          when pause_getII3771 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1414\ := \$arr1452_value\;
            if \$1414_lock\(0) = '1' then
              \state\ <= get_wait3769;
            else
              \$1398\ := \$1414\;
              \$v3768\ := \$arr1452_ptr_take\;
              if \$v3768\(0) = '1' then
                \state\ <= q_wait3767;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3765;
              end if;
            end if;
          when pause_getII3779 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1430\ := \$arr1451_value\;
            \$1428\ := \$1430\(36 to 71);
            \$v3776\ := \$1428\;
            \$v3777\ := \$v3776\(0 to 3);
            \$v3775\ := \$v3776\(4 to 35);
            case \$v3777\ is
            when "0010" =>
              \$1397\ := eclat_true;
              \$v3774\ := \$1397\;
              if \$v3774\(0) = '1' then
                \$v3745\ := \$arr1452_ptr_take\;
                if \$v3745\(0) = '1' then
                  \state\ <= q_wait3744;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3742;
                end if;
              else
                \$v3773\ := \$arr1452_ptr_take\;
                if \$v3773\(0) = '1' then
                  \state\ <= q_wait3772;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3770;
                end if;
              end if;
            when others =>
              \$1397\ := eclat_false;
              \$v3774\ := \$1397\;
              if \$v3774\(0) = '1' then
                \$v3745\ := \$arr1452_ptr_take\;
                if \$v3745\(0) = '1' then
                  \state\ <= q_wait3744;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3742;
                end if;
              else
                \$v3773\ := \$arr1452_ptr_take\;
                if \$v3773\(0) = '1' then
                  \state\ <= q_wait3772;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3770;
                end if;
              end if;
            end case;
          when pause_getII3784 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1435\ := \$arr1452_value\;
            if \$1435_lock\(0) = '1' then
              \state\ <= get_wait3782;
            else
              \$1434\ := \$1435\;
              \$v3781\ := \$arr1451_ptr_take\;
              if \$v3781\(0) = '1' then
                \state\ <= q_wait3780;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1434\));
                \state\ <= pause_getI3778;
              end if;
            end if;
          when pause_getII3788 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1436\ := \$arr1451_value\;
            \$1396_x\ := \$1436\(0 to 35);
            \$v3786\ := \$arr1452_ptr_take\;
            if \$v3786\(0) = '1' then
              \state\ <= q_wait3785;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3783;
            end if;
          when pause_getII3793 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1441\ := \$arr1452_value\;
            if \$1441_lock\(0) = '1' then
              \state\ <= get_wait3791;
            else
              \$1440\ := \$1441\;
              \$v3790\ := \$arr1451_ptr_take\;
              if \$v3790\(0) = '1' then
                \state\ <= q_wait3789;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1440\));
                \state\ <= pause_getI3787;
              end if;
            end if;
          when pause_getII3802 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1468\ := \$arr1451_value\;
            \$1463\ := \$1468\(36 to 71);
            \$v3799\ := \$1463\;
            \$v3800\ := \$v3799\(0 to 3);
            \$v3798\ := \$v3799\(4 to 35);
            case \$v3800\ is
            when "0010" =>
              \$1464_i\ := \$v3798\(0 to 31);
              \$1462\ := \$1464_i\;
              if \$1461_lock\(0) = '1' then
                \state\ <= get_wait3796;
              else
                \$1461_lock\ := eclat_true;
                \state\ <= get_pause3797;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811444\;
            end case;
          when pause_getII3807 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1473\ := \$arr1452_value\;
            if \$1473_lock\(0) = '1' then
              \state\ <= get_wait3805;
            else
              \$1472\ := \$1473\;
              \$v3804\ := \$arr1451_ptr_take\;
              if \$v3804\(0) = '1' then
                \state\ <= q_wait3803;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1472\));
                \state\ <= pause_getI3801;
              end if;
            end if;
          when pause_getII3811 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3809\ := \$arr1452_ptr_take\;
            if \$v3809\(0) = '1' then
              \state\ <= q_wait3808;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3806;
            end if;
          when pause_getII3820 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1448\ := \$arr1451_value\;
            \$1447\ := \$1448\(72 to 107);
            \$v3818\ := "00000000000000000000000000000000";
            \$1445\ := "0000" & \$v3818\ & \$1446\ & \$1447\;
            \$v3817\ := \$arr1451_ptr_take\;
            if \$v3817\(0) = '1' then
              \state\ <= q_wait3816;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1444\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1445\;
              \state\ <= pause_setI3814;
            end if;
          when pause_getII3825 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1453\ := \$arr1452_value\;
            if \$1453_lock\(0) = '1' then
              \state\ <= get_wait3823;
            else
              \$1452\ := \$1453\;
              \$v3822\ := \$arr1451_ptr_take\;
              if \$v3822\(0) = '1' then
                \state\ <= q_wait3821;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1452\));
                \state\ <= pause_getI3819;
              end if;
            end if;
          when pause_getII3829 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1454\ := \$arr1451_value\;
            \$1446\ := \$1454\(36 to 71);
            \$v3827\ := \$arr1452_ptr_take\;
            if \$v3827\(0) = '1' then
              \state\ <= q_wait3826;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3824;
            end if;
          when pause_getII3834 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1459\ := \$arr1452_value\;
            if \$1459_lock\(0) = '1' then
              \state\ <= get_wait3832;
            else
              \$1458\ := \$1459\;
              \$v3831\ := \$arr1451_ptr_take\;
              if \$v3831\(0) = '1' then
                \state\ <= q_wait3830;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1458\));
                \state\ <= pause_getI3828;
              end if;
            end if;
          when pause_getII3839 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1460\ := \$arr1452_value\;
            if \$1460_lock\(0) = '1' then
              \state\ <= get_wait3837;
            else
              \$1444\ := \$1460\;
              \$v3836\ := \$arr1452_ptr_take\;
              if \$v3836\(0) = '1' then
                \state\ <= q_wait3835;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3833;
              end if;
            end if;
          when pause_getII3847 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1476\ := \$arr1451_value\;
            \$1474\ := \$1476\(36 to 71);
            \$v3844\ := \$1474\;
            \$v3845\ := \$v3844\(0 to 3);
            \$v3843\ := \$v3844\(4 to 35);
            case \$v3845\ is
            when "0010" =>
              \$1443\ := eclat_true;
              \$v3842\ := \$1443\;
              if \$v3842\(0) = '1' then
                \$v3813\ := \$arr1452_ptr_take\;
                if \$v3813\(0) = '1' then
                  \state\ <= q_wait3812;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3810;
                end if;
              else
                \$v3841\ := \$arr1452_ptr_take\;
                if \$v3841\(0) = '1' then
                  \state\ <= q_wait3840;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3838;
                end if;
              end if;
            when others =>
              \$1443\ := eclat_false;
              \$v3842\ := \$1443\;
              if \$v3842\(0) = '1' then
                \$v3813\ := \$arr1452_ptr_take\;
                if \$v3813\(0) = '1' then
                  \state\ <= q_wait3812;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3810;
                end if;
              else
                \$v3841\ := \$arr1452_ptr_take\;
                if \$v3841\(0) = '1' then
                  \state\ <= q_wait3840;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3838;
                end if;
              end if;
            end case;
          when pause_getII3852 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1481\ := \$arr1452_value\;
            if \$1481_lock\(0) = '1' then
              \state\ <= get_wait3850;
            else
              \$1480\ := \$1481\;
              \$v3849\ := \$arr1451_ptr_take\;
              if \$v3849\(0) = '1' then
                \state\ <= q_wait3848;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1480\));
                \state\ <= pause_getI3846;
              end if;
            end if;
          when pause_getII3856 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1482\ := \$arr1451_value\;
            \$1442_x\ := \$1482\(0 to 35);
            \$v3854\ := \$arr1452_ptr_take\;
            if \$v3854\(0) = '1' then
              \state\ <= q_wait3853;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3851;
            end if;
          when pause_getII3861 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1487\ := \$arr1452_value\;
            if \$1487_lock\(0) = '1' then
              \state\ <= get_wait3859;
            else
              \$1486\ := \$1487\;
              \$v3858\ := \$arr1451_ptr_take\;
              if \$v3858\(0) = '1' then
                \state\ <= q_wait3857;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1486\));
                \state\ <= pause_getI3855;
              end if;
            end if;
          when pause_getII3872 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1497\ := \$arr1452_value\;
            if \$1497_lock\(0) = '1' then
              \state\ <= get_wait3870;
            else
              \$1496\ := \$1497\;
              \$1495\ := \$1496\ & "00000000000000000000000000000001";
              \$1494\ := eclat_sub(\$1495\);
              if \$1493_lock\(0) = '1' then
                \state\ <= get_wait3868;
              else
                \$1493_lock\ := eclat_true;
                \state\ <= get_pause3869;
              end if;
            end if;
          when pause_getII3876 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3874\ := \$arr1452_ptr_take\;
            if \$v3874\(0) = '1' then
              \state\ <= q_wait3873;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3871;
            end if;
          when pause_getII3888 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1492_lock\(0) = '1' then
              \state\ <= get_wait3885;
            else
              \$1492_lock\ := eclat_true;
              \state\ <= get_pause3886;
            end if;
          when pause_getII3900 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1498\ := \$arr1452_value\;
            if \$1498_lock\(0) = '1' then
              \state\ <= get_wait3898;
            else
              \$1488_i\ := \$1498\;
              \$v3897\ := eclat_gt(\$1488_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v3897\(0) = '1' then
                \$v3896\ := eclat_eq(\$1488_i\ & X"000" & X"15f90");
                if \$v3896\(0) = '1' then
                  \$v3884\ := \$arr1451_ptr_take\;
                  if \$v3884\(0) = '1' then
                    \state\ <= q_wait3883;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3879\ := "00000000000000000000000000000000";
                    \$v3880\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$76_result\ & "0001" & \$v3879\ & "0001" & \$v3880\;
                    \state\ <= pause_setI3881;
                  end if;
                else
                  \$v3895\ := \$arr1451_ptr_take\;
                  if \$v3895\(0) = '1' then
                    \state\ <= q_wait3894;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$v3891\ := "00000000000000000000000000000000";
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$76_result\ & "0010" & \$1488_i\ & "0001" & \$v3891\;
                    \state\ <= pause_setI3892;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811445\;
              end if;
            end if;
          when pause_getII3909 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1525\ := \$arr1451_value\;
            \$1520\ := \$1525\(36 to 71);
            \$v3906\ := \$1520\;
            \$v3907\ := \$v3906\(0 to 3);
            \$v3905\ := \$v3906\(4 to 35);
            case \$v3907\ is
            when "0010" =>
              \$1521_i\ := \$v3905\(0 to 31);
              \$1519\ := \$1521_i\;
              if \$1518_lock\(0) = '1' then
                \state\ <= get_wait3903;
              else
                \$1518_lock\ := eclat_true;
                \state\ <= get_pause3904;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811446\;
            end case;
          when pause_getII3914 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1530\ := \$arr1452_value\;
            if \$1530_lock\(0) = '1' then
              \state\ <= get_wait3912;
            else
              \$1529\ := \$1530\;
              \$v3911\ := \$arr1451_ptr_take\;
              if \$v3911\(0) = '1' then
                \state\ <= q_wait3910;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1529\));
                \state\ <= pause_getI3908;
              end if;
            end if;
          when pause_getII3918 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v3916\ := \$arr1452_ptr_take\;
            if \$v3916\(0) = '1' then
              \state\ <= q_wait3915;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3913;
            end if;
          when pause_getII3927 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1505\ := \$arr1451_value\;
            \$1504\ := \$1505\(72 to 107);
            \$v3925\ := "00000000000000000000000000000000";
            \$1502\ := "0000" & \$v3925\ & \$1503\ & \$1504\;
            \$v3924\ := \$arr1451_ptr_take\;
            if \$v3924\(0) = '1' then
              \state\ <= q_wait3923;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1501\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1502\;
              \state\ <= pause_setI3921;
            end if;
          when pause_getII3932 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1510\ := \$arr1452_value\;
            if \$1510_lock\(0) = '1' then
              \state\ <= get_wait3930;
            else
              \$1509\ := \$1510\;
              \$v3929\ := \$arr1451_ptr_take\;
              if \$v3929\(0) = '1' then
                \state\ <= q_wait3928;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1509\));
                \state\ <= pause_getI3926;
              end if;
            end if;
          when pause_getII3936 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1511\ := \$arr1451_value\;
            \$1503\ := \$1511\(36 to 71);
            \$v3934\ := \$arr1452_ptr_take\;
            if \$v3934\(0) = '1' then
              \state\ <= q_wait3933;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3931;
            end if;
          when pause_getII3941 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1516\ := \$arr1452_value\;
            if \$1516_lock\(0) = '1' then
              \state\ <= get_wait3939;
            else
              \$1515\ := \$1516\;
              \$v3938\ := \$arr1451_ptr_take\;
              if \$v3938\(0) = '1' then
                \state\ <= q_wait3937;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1515\));
                \state\ <= pause_getI3935;
              end if;
            end if;
          when pause_getII3946 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1517\ := \$arr1452_value\;
            if \$1517_lock\(0) = '1' then
              \state\ <= get_wait3944;
            else
              \$1501\ := \$1517\;
              \$v3943\ := \$arr1452_ptr_take\;
              if \$v3943\(0) = '1' then
                \state\ <= q_wait3942;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3940;
              end if;
            end if;
          when pause_getII3954 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1533\ := \$arr1451_value\;
            \$1531\ := \$1533\(36 to 71);
            \$v3951\ := \$1531\;
            \$v3952\ := \$v3951\(0 to 3);
            \$v3950\ := \$v3951\(4 to 35);
            case \$v3952\ is
            when "0010" =>
              \$1500\ := eclat_true;
              \$v3949\ := \$1500\;
              if \$v3949\(0) = '1' then
                \$v3920\ := \$arr1452_ptr_take\;
                if \$v3920\(0) = '1' then
                  \state\ <= q_wait3919;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3917;
                end if;
              else
                \$v3948\ := \$arr1452_ptr_take\;
                if \$v3948\(0) = '1' then
                  \state\ <= q_wait3947;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3945;
                end if;
              end if;
            when others =>
              \$1500\ := eclat_false;
              \$v3949\ := \$1500\;
              if \$v3949\(0) = '1' then
                \$v3920\ := \$arr1452_ptr_take\;
                if \$v3920\(0) = '1' then
                  \state\ <= q_wait3919;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3917;
                end if;
              else
                \$v3948\ := \$arr1452_ptr_take\;
                if \$v3948\(0) = '1' then
                  \state\ <= q_wait3947;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI3945;
                end if;
              end if;
            end case;
          when pause_getII3959 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1538\ := \$arr1452_value\;
            if \$1538_lock\(0) = '1' then
              \state\ <= get_wait3957;
            else
              \$1537\ := \$1538\;
              \$v3956\ := \$arr1451_ptr_take\;
              if \$v3956\(0) = '1' then
                \state\ <= q_wait3955;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1537\));
                \state\ <= pause_getI3953;
              end if;
            end if;
          when pause_getII3963 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1539\ := \$arr1451_value\;
            \$1499_x\ := \$1539\(0 to 35);
            \$v3961\ := \$arr1452_ptr_take\;
            if \$v3961\(0) = '1' then
              \state\ <= q_wait3960;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3958;
            end if;
          when pause_getII3968 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1544\ := \$arr1452_value\;
            if \$1544_lock\(0) = '1' then
              \state\ <= get_wait3966;
            else
              \$1543\ := \$1544\;
              \$v3965\ := \$arr1451_ptr_take\;
              if \$v3965\(0) = '1' then
                \state\ <= q_wait3964;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1543\));
                \state\ <= pause_getI3962;
              end if;
            end if;
          when pause_getII3978 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1550_lock\(0) = '1' then
              \state\ <= get_wait3975;
            else
              \$1550_lock\ := eclat_true;
              \state\ <= get_pause3976;
            end if;
          when pause_getII3988 =>
            \$arr1452_ptr_take\(0) := '0';
            if \$1549_lock\(0) = '1' then
              \state\ <= get_wait3985;
            else
              \$1549_lock\ := eclat_true;
              \state\ <= get_pause3986;
            end if;
          when pause_getII4005 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1551\ := \$arr1452_value\;
            if \$1551_lock\(0) = '1' then
              \state\ <= get_wait4003;
            else
              \$1545_i\ := \$1551\;
              \$v4002\ := eclat_gt(\$1545_i\ & eclat_sub(eclat_div(X"000" & X"15f90" & "00000000000000000000000000000010") & "00000000000000000000000000000001"));
              if \$v4002\(0) = '1' then
                \$v4001\ := eclat_eq(\$1545_i\ & X"000" & X"15f90");
                if \$v4001\(0) = '1' then
                  \$v3984\ := \$arr1451_ptr_take\;
                  if \$v3984\(0) = '1' then
                    \state\ <= q_wait3983;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
                    \state\ <= pause_setI3981;
                  end if;
                else
                  \$v4000\ := \$arr1451_ptr_take\;
                  if \$v4000\(0) = '1' then
                    \state\ <= q_wait3999;
                  else
                    \$arr1451_ptr_take\(0) := '1';
                    \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
                    \$arr1451_write_request\ <= '1';
                    \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
                    \state\ <= pause_setI3997;
                  end if;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("stack overflow"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811447\;
              end if;
            end if;
          when pause_getII4014 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1578\ := \$arr1451_value\;
            \$1573\ := \$1578\(36 to 71);
            \$v4011\ := \$1573\;
            \$v4012\ := \$v4011\(0 to 3);
            \$v4010\ := \$v4011\(4 to 35);
            case \$v4012\ is
            when "0010" =>
              \$1574_i\ := \$v4010\(0 to 31);
              \$1572\ := \$1574_i\;
              if \$1571_lock\(0) = '1' then
                \state\ <= get_wait4008;
              else
                \$1571_lock\ := eclat_true;
                \state\ <= get_pause4009;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811448\;
            end case;
          when pause_getII4019 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1583\ := \$arr1452_value\;
            if \$1583_lock\(0) = '1' then
              \state\ <= get_wait4017;
            else
              \$1582\ := \$1583\;
              \$v4016\ := \$arr1451_ptr_take\;
              if \$v4016\(0) = '1' then
                \state\ <= q_wait4015;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1582\));
                \state\ <= pause_getI4013;
              end if;
            end if;
          when pause_getII4023 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4021\ := \$arr1452_ptr_take\;
            if \$v4021\(0) = '1' then
              \state\ <= q_wait4020;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4018;
            end if;
          when pause_getII4032 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1558\ := \$arr1451_value\;
            \$1557\ := \$1558\(72 to 107);
            \$v4030\ := "00000000000000000000000000000000";
            \$1555\ := "0000" & \$v4030\ & \$1556\ & \$1557\;
            \$v4029\ := \$arr1451_ptr_take\;
            if \$v4029\(0) = '1' then
              \state\ <= q_wait4028;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1554\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1555\;
              \state\ <= pause_setI4026;
            end if;
          when pause_getII4037 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1563\ := \$arr1452_value\;
            if \$1563_lock\(0) = '1' then
              \state\ <= get_wait4035;
            else
              \$1562\ := \$1563\;
              \$v4034\ := \$arr1451_ptr_take\;
              if \$v4034\(0) = '1' then
                \state\ <= q_wait4033;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1562\));
                \state\ <= pause_getI4031;
              end if;
            end if;
          when pause_getII4041 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1564\ := \$arr1451_value\;
            \$1556\ := \$1564\(36 to 71);
            \$v4039\ := \$arr1452_ptr_take\;
            if \$v4039\(0) = '1' then
              \state\ <= q_wait4038;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4036;
            end if;
          when pause_getII4046 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1569\ := \$arr1452_value\;
            if \$1569_lock\(0) = '1' then
              \state\ <= get_wait4044;
            else
              \$1568\ := \$1569\;
              \$v4043\ := \$arr1451_ptr_take\;
              if \$v4043\(0) = '1' then
                \state\ <= q_wait4042;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1568\));
                \state\ <= pause_getI4040;
              end if;
            end if;
          when pause_getII4051 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1570\ := \$arr1452_value\;
            if \$1570_lock\(0) = '1' then
              \state\ <= get_wait4049;
            else
              \$1554\ := \$1570\;
              \$v4048\ := \$arr1452_ptr_take\;
              if \$v4048\(0) = '1' then
                \state\ <= q_wait4047;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4045;
              end if;
            end if;
          when pause_getII4059 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1586\ := \$arr1451_value\;
            \$1584\ := \$1586\(36 to 71);
            \$v4056\ := \$1584\;
            \$v4057\ := \$v4056\(0 to 3);
            \$v4055\ := \$v4056\(4 to 35);
            case \$v4057\ is
            when "0010" =>
              \$1553\ := eclat_true;
              \$v4054\ := \$1553\;
              if \$v4054\(0) = '1' then
                \$v4025\ := \$arr1452_ptr_take\;
                if \$v4025\(0) = '1' then
                  \state\ <= q_wait4024;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4022;
                end if;
              else
                \$v4053\ := \$arr1452_ptr_take\;
                if \$v4053\(0) = '1' then
                  \state\ <= q_wait4052;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4050;
                end if;
              end if;
            when others =>
              \$1553\ := eclat_false;
              \$v4054\ := \$1553\;
              if \$v4054\(0) = '1' then
                \$v4025\ := \$arr1452_ptr_take\;
                if \$v4025\(0) = '1' then
                  \state\ <= q_wait4024;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4022;
                end if;
              else
                \$v4053\ := \$arr1452_ptr_take\;
                if \$v4053\(0) = '1' then
                  \state\ <= q_wait4052;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4050;
                end if;
              end if;
            end case;
          when pause_getII4064 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1591\ := \$arr1452_value\;
            if \$1591_lock\(0) = '1' then
              \state\ <= get_wait4062;
            else
              \$1590\ := \$1591\;
              \$v4061\ := \$arr1451_ptr_take\;
              if \$v4061\(0) = '1' then
                \state\ <= q_wait4060;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1590\));
                \state\ <= pause_getI4058;
              end if;
            end if;
          when pause_getII4068 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1592\ := \$arr1451_value\;
            \$1552_x\ := \$1592\(0 to 35);
            \$v4066\ := \$arr1452_ptr_take\;
            if \$v4066\(0) = '1' then
              \state\ <= q_wait4065;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4063;
            end if;
          when pause_getII4073 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1597\ := \$arr1452_value\;
            if \$1597_lock\(0) = '1' then
              \state\ <= get_wait4071;
            else
              \$1596\ := \$1597\;
              \$v4070\ := \$arr1451_ptr_take\;
              if \$v4070\(0) = '1' then
                \state\ <= q_wait4069;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1596\));
                \state\ <= pause_getI4067;
              end if;
            end if;
          when pause_getII4082 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1624\ := \$arr1451_value\;
            \$1619\ := \$1624\(36 to 71);
            \$v4079\ := \$1619\;
            \$v4080\ := \$v4079\(0 to 3);
            \$v4078\ := \$v4079\(4 to 35);
            case \$v4080\ is
            when "0010" =>
              \$1620_i\ := \$v4078\(0 to 31);
              \$1618\ := \$1620_i\;
              if \$1617_lock\(0) = '1' then
                \state\ <= get_wait4076;
              else
                \$1617_lock\ := eclat_true;
                \state\ <= get_pause4077;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811449\;
            end case;
          when pause_getII4087 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1629\ := \$arr1452_value\;
            if \$1629_lock\(0) = '1' then
              \state\ <= get_wait4085;
            else
              \$1628\ := \$1629\;
              \$v4084\ := \$arr1451_ptr_take\;
              if \$v4084\(0) = '1' then
                \state\ <= q_wait4083;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1628\));
                \state\ <= pause_getI4081;
              end if;
            end if;
          when pause_getII4091 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4089\ := \$arr1452_ptr_take\;
            if \$v4089\(0) = '1' then
              \state\ <= q_wait4088;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4086;
            end if;
          when pause_getII4100 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1604\ := \$arr1451_value\;
            \$1603\ := \$1604\(72 to 107);
            \$v4098\ := "00000000000000000000000000000000";
            \$1601\ := "0000" & \$v4098\ & \$1602\ & \$1603\;
            \$v4097\ := \$arr1451_ptr_take\;
            if \$v4097\(0) = '1' then
              \state\ <= q_wait4096;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1600\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1601\;
              \state\ <= pause_setI4094;
            end if;
          when pause_getII4105 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1609\ := \$arr1452_value\;
            if \$1609_lock\(0) = '1' then
              \state\ <= get_wait4103;
            else
              \$1608\ := \$1609\;
              \$v4102\ := \$arr1451_ptr_take\;
              if \$v4102\(0) = '1' then
                \state\ <= q_wait4101;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1608\));
                \state\ <= pause_getI4099;
              end if;
            end if;
          when pause_getII4109 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1610\ := \$arr1451_value\;
            \$1602\ := \$1610\(36 to 71);
            \$v4107\ := \$arr1452_ptr_take\;
            if \$v4107\(0) = '1' then
              \state\ <= q_wait4106;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4104;
            end if;
          when pause_getII4114 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1615\ := \$arr1452_value\;
            if \$1615_lock\(0) = '1' then
              \state\ <= get_wait4112;
            else
              \$1614\ := \$1615\;
              \$v4111\ := \$arr1451_ptr_take\;
              if \$v4111\(0) = '1' then
                \state\ <= q_wait4110;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1614\));
                \state\ <= pause_getI4108;
              end if;
            end if;
          when pause_getII4119 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1616\ := \$arr1452_value\;
            if \$1616_lock\(0) = '1' then
              \state\ <= get_wait4117;
            else
              \$1600\ := \$1616\;
              \$v4116\ := \$arr1452_ptr_take\;
              if \$v4116\(0) = '1' then
                \state\ <= q_wait4115;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4113;
              end if;
            end if;
          when pause_getII4127 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1632\ := \$arr1451_value\;
            \$1630\ := \$1632\(36 to 71);
            \$v4124\ := \$1630\;
            \$v4125\ := \$v4124\(0 to 3);
            \$v4123\ := \$v4124\(4 to 35);
            case \$v4125\ is
            when "0010" =>
              \$1599\ := eclat_true;
              \$v4122\ := \$1599\;
              if \$v4122\(0) = '1' then
                \$v4093\ := \$arr1452_ptr_take\;
                if \$v4093\(0) = '1' then
                  \state\ <= q_wait4092;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4090;
                end if;
              else
                \$v4121\ := \$arr1452_ptr_take\;
                if \$v4121\(0) = '1' then
                  \state\ <= q_wait4120;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4118;
                end if;
              end if;
            when others =>
              \$1599\ := eclat_false;
              \$v4122\ := \$1599\;
              if \$v4122\(0) = '1' then
                \$v4093\ := \$arr1452_ptr_take\;
                if \$v4093\(0) = '1' then
                  \state\ <= q_wait4092;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4090;
                end if;
              else
                \$v4121\ := \$arr1452_ptr_take\;
                if \$v4121\(0) = '1' then
                  \state\ <= q_wait4120;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4118;
                end if;
              end if;
            end case;
          when pause_getII4132 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1637\ := \$arr1452_value\;
            if \$1637_lock\(0) = '1' then
              \state\ <= get_wait4130;
            else
              \$1636\ := \$1637\;
              \$v4129\ := \$arr1451_ptr_take\;
              if \$v4129\(0) = '1' then
                \state\ <= q_wait4128;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1636\));
                \state\ <= pause_getI4126;
              end if;
            end if;
          when pause_getII4136 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1638\ := \$arr1451_value\;
            \$1598_x\ := \$1638\(0 to 35);
            \$v4134\ := \$arr1452_ptr_take\;
            if \$v4134\(0) = '1' then
              \state\ <= q_wait4133;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4131;
            end if;
          when pause_getII4141 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1643\ := \$arr1452_value\;
            if \$1643_lock\(0) = '1' then
              \state\ <= get_wait4139;
            else
              \$1642\ := \$1643\;
              \$v4138\ := \$arr1451_ptr_take\;
              if \$v4138\(0) = '1' then
                \state\ <= q_wait4137;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1642\));
                \state\ <= pause_getI4135;
              end if;
            end if;
          when pause_getII4150 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1670\ := \$arr1451_value\;
            \$1665\ := \$1670\(36 to 71);
            \$v4147\ := \$1665\;
            \$v4148\ := \$v4147\(0 to 3);
            \$v4146\ := \$v4147\(4 to 35);
            case \$v4148\ is
            when "0010" =>
              \$1666_i\ := \$v4146\(0 to 31);
              \$1664\ := \$1666_i\;
              if \$1663_lock\(0) = '1' then
                \state\ <= get_wait4144;
              else
                \$1663_lock\ := eclat_true;
                \state\ <= get_pause4145;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811450\;
            end case;
          when pause_getII4155 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1675\ := \$arr1452_value\;
            if \$1675_lock\(0) = '1' then
              \state\ <= get_wait4153;
            else
              \$1674\ := \$1675\;
              \$v4152\ := \$arr1451_ptr_take\;
              if \$v4152\(0) = '1' then
                \state\ <= q_wait4151;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1674\));
                \state\ <= pause_getI4149;
              end if;
            end if;
          when pause_getII4159 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4157\ := \$arr1452_ptr_take\;
            if \$v4157\(0) = '1' then
              \state\ <= q_wait4156;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4154;
            end if;
          when pause_getII4168 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1650\ := \$arr1451_value\;
            \$1649\ := \$1650\(72 to 107);
            \$v4166\ := "00000000000000000000000000000000";
            \$1647\ := "0000" & \$v4166\ & \$1648\ & \$1649\;
            \$v4165\ := \$arr1451_ptr_take\;
            if \$v4165\(0) = '1' then
              \state\ <= q_wait4164;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1646\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1647\;
              \state\ <= pause_setI4162;
            end if;
          when pause_getII4173 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1655\ := \$arr1452_value\;
            if \$1655_lock\(0) = '1' then
              \state\ <= get_wait4171;
            else
              \$1654\ := \$1655\;
              \$v4170\ := \$arr1451_ptr_take\;
              if \$v4170\(0) = '1' then
                \state\ <= q_wait4169;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1654\));
                \state\ <= pause_getI4167;
              end if;
            end if;
          when pause_getII4177 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1656\ := \$arr1451_value\;
            \$1648\ := \$1656\(36 to 71);
            \$v4175\ := \$arr1452_ptr_take\;
            if \$v4175\(0) = '1' then
              \state\ <= q_wait4174;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4172;
            end if;
          when pause_getII4182 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1661\ := \$arr1452_value\;
            if \$1661_lock\(0) = '1' then
              \state\ <= get_wait4180;
            else
              \$1660\ := \$1661\;
              \$v4179\ := \$arr1451_ptr_take\;
              if \$v4179\(0) = '1' then
                \state\ <= q_wait4178;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1660\));
                \state\ <= pause_getI4176;
              end if;
            end if;
          when pause_getII4187 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1662\ := \$arr1452_value\;
            if \$1662_lock\(0) = '1' then
              \state\ <= get_wait4185;
            else
              \$1646\ := \$1662\;
              \$v4184\ := \$arr1452_ptr_take\;
              if \$v4184\(0) = '1' then
                \state\ <= q_wait4183;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI4181;
              end if;
            end if;
          when pause_getII4195 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1678\ := \$arr1451_value\;
            \$1676\ := \$1678\(36 to 71);
            \$v4192\ := \$1676\;
            \$v4193\ := \$v4192\(0 to 3);
            \$v4191\ := \$v4192\(4 to 35);
            case \$v4193\ is
            when "0010" =>
              \$1645\ := eclat_true;
              \$v4190\ := \$1645\;
              if \$v4190\(0) = '1' then
                \$v4161\ := \$arr1452_ptr_take\;
                if \$v4161\(0) = '1' then
                  \state\ <= q_wait4160;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4158;
                end if;
              else
                \$v4189\ := \$arr1452_ptr_take\;
                if \$v4189\(0) = '1' then
                  \state\ <= q_wait4188;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4186;
                end if;
              end if;
            when others =>
              \$1645\ := eclat_false;
              \$v4190\ := \$1645\;
              if \$v4190\(0) = '1' then
                \$v4161\ := \$arr1452_ptr_take\;
                if \$v4161\(0) = '1' then
                  \state\ <= q_wait4160;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4158;
                end if;
              else
                \$v4189\ := \$arr1452_ptr_take\;
                if \$v4189\(0) = '1' then
                  \state\ <= q_wait4188;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI4186;
                end if;
              end if;
            end case;
          when pause_getII4200 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1683\ := \$arr1452_value\;
            if \$1683_lock\(0) = '1' then
              \state\ <= get_wait4198;
            else
              \$1682\ := \$1683\;
              \$v4197\ := \$arr1451_ptr_take\;
              if \$v4197\(0) = '1' then
                \state\ <= q_wait4196;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1682\));
                \state\ <= pause_getI4194;
              end if;
            end if;
          when pause_getII4204 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1684\ := \$arr1451_value\;
            \$1644_x\ := \$1684\(0 to 35);
            \$v4202\ := \$arr1452_ptr_take\;
            if \$v4202\(0) = '1' then
              \state\ <= q_wait4201;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4199;
            end if;
          when pause_getII4209 =>
            \$arr1452_ptr_take\(0) := '0';
            \$1689\ := \$arr1452_value\;
            if \$1689_lock\(0) = '1' then
              \state\ <= get_wait4207;
            else
              \$1688\ := \$1689\;
              \$v4206\ := \$arr1451_ptr_take\;
              if \$v4206\(0) = '1' then
                \state\ <= q_wait4205;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1688\));
                \state\ <= pause_getI4203;
              end if;
            end if;
          when pause_getII4213 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v18\ := \$arr1451_value\;
            \$v4211\ := \$arr1452_ptr_take\;
            if \$v4211\(0) = '1' then
              \state\ <= q_wait4210;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4208;
            end if;
          when pause_getII4218 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v16\ := \$arr1452_value\;
            if \$v16_lock\(0) = '1' then
              \state\ <= get_wait4216;
            else
              \$v17\ := \$v16\;
              \$v4215\ := \$arr1451_ptr_take\;
              if \$v4215\(0) = '1' then
                \state\ <= q_wait4214;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$v17\));
                \state\ <= pause_getI4212;
              end if;
            end if;
          when pause_setI1457 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII1458;
          when pause_setI1474 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1475;
          when pause_setI1485 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1486;
          when pause_setI1521 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1522;
          when pause_setI1589 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1590;
          when pause_setI1639 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII1640;
          when pause_setI1656 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1657;
          when pause_setI1667 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1668;
          when pause_setI1703 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1704;
          when pause_setI1771 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1772;
          when pause_setI1821 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII1822;
          when pause_setI1838 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1839;
          when pause_setI1849 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1850;
          when pause_setI1885 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1886;
          when pause_setI1953 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII1954;
          when pause_setI2003 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2004;
          when pause_setI2020 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2021;
          when pause_setI2031 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2032;
          when pause_setI2067 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2068;
          when pause_setI2135 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2136;
          when pause_setI2185 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2186;
          when pause_setI2201 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2202;
          when pause_setI2213 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2214;
          when pause_setI2223 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2224;
          when pause_setI2258 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2259;
          when pause_setI2326 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2327;
          when pause_setI2376 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2377;
          when pause_setI2392 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2393;
          when pause_setI2404 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2405;
          when pause_setI2414 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2415;
          when pause_setI2452 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2453;
          when pause_setI2520 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2521;
          when pause_setI2570 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2571;
          when pause_setI2580 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2581;
          when pause_setI2592 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2593;
          when pause_setI2596 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2597;
          when pause_setI2632 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2633;
          when pause_setI2700 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2701;
          when pause_setI2750 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2751;
          when pause_setI2760 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2761;
          when pause_setI2772 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2773;
          when pause_setI2776 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2777;
          when pause_setI2812 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2813;
          when pause_setI2880 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2881;
          when pause_setI2930 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII2931;
          when pause_setI2940 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2941;
          when pause_setI2952 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2953;
          when pause_setI2956 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2957;
          when pause_setI2992 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII2993;
          when pause_setI3060 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3061;
          when pause_setI3110 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3111;
          when pause_setI3127 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3128;
          when pause_setI3138 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3139;
          when pause_setI3174 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3175;
          when pause_setI3224 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3225;
          when pause_setI3241 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3242;
          when pause_setI3252 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3253;
          when pause_setI3288 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3289;
          when pause_setI3338 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3339;
          when pause_setI3355 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3356;
          when pause_setI3366 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3367;
          when pause_setI3402 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3403;
          when pause_setI3452 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3453;
          when pause_setI3462 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3463;
          when pause_setI3474 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3475;
          when pause_setI3478 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3479;
          when pause_setI3516 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3517;
          when pause_setI3566 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3567;
          when pause_setI3577 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3578;
          when pause_setI3589 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3590;
          when pause_setI3594 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3595;
          when pause_setI3639 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3640;
          when pause_setI3689 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3690;
          when pause_setI3706 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3707;
          when pause_setI3717 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3718;
          when pause_setI3746 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3747;
          when pause_setI3814 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3815;
          when pause_setI3864 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3865;
          when pause_setI3881 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3882;
          when pause_setI3892 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3893;
          when pause_setI3921 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3922;
          when pause_setI3971 =>
            \$arr1453_write_request\ <= '0';
            \state\ <= pause_setII3972;
          when pause_setI3981 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3982;
          when pause_setI3993 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3994;
          when pause_setI3997 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII3998;
          when pause_setI4026 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII4027;
          when pause_setI4094 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII4095;
          when pause_setI4162 =>
            \$arr1451_write_request\ <= '0';
            \state\ <= pause_setII4163;
          when pause_setI4221 =>
            \$arr1452_write_request\ <= '0';
            \state\ <= pause_setII4222;
          when pause_setI4225 =>
            \$arr1452_write_request\ <= '0';
            \state\ <= pause_setII4226;
          when pause_setI4229 =>
            \$arr1452_write_request\ <= '0';
            \state\ <= pause_setII4230;
          when pause_setI4233 =>
            \$arr1452_write_request\ <= '0';
            \state\ <= pause_setII4234;
          when pause_setI4237 =>
            \$arr1452_write_request\ <= '0';
            \state\ <= pause_setII4238;
          when pause_setII1458 =>
            \$arr1453_ptr_take\(0) := '0';
            result1454 := eclat_unit;
            eclat_print_string(of_string("Test"));
            
            rdy1455 := eclat_true;
            \state\ <= compute1456;
          when pause_setII1475 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1471\ := \$arr1452_ptr_take\;
            if \$v1471\(0) = '1' then
              \state\ <= q_wait1470;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1468;
            end if;
          when pause_setII1486 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1483\ := \$arr1452_ptr_take\;
            if \$v1483\(0) = '1' then
              \state\ <= q_wait1482;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1480;
            end if;
          when pause_setII1522 =>
            \$arr1451_ptr_take\(0) := '0';
            \$70_y\ := \$84_x\;
            \$v1501\ := \$70_y\;
            \$v1502\ := \$v1501\(0 to 3);
            \$v1496\ := \$v1501\(4 to 35);
            case \$v1502\ is
            when "0001" =>
              a := \$v1496\(0 to 31);
              \$v1499\ := \$69_x\;
              \$v1500\ := \$v1499\(0 to 3);
              \$v1497\ := \$v1499\(4 to 35);
              case \$v1500\ is
              when "0001" =>
                b := \$v1497\(0 to 31);
                \$v1498\ := eclat_div(a & b);
                \$71_result_after_f\ := "0001" & \$v1498\;
                \$v1495\ := \$arr1452_ptr_take\;
                if \$v1495\(0) = '1' then
                  \state\ <= q_wait1494;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1492;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("* quotient arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811390\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("* quotient arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811389\;
            end case;
          when pause_setII1590 =>
            \$arr1451_ptr_take\(0) := '0';
            \$69_x\ := \$161_x\;
            \$v1570\ := \$arr1452_ptr_take\;
            if \$v1570\(0) = '1' then
              \state\ <= q_wait1569;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1567;
            end if;
          when pause_setII1640 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v1638\ := \$arr1452_ptr_take\;
            if \$v1638\(0) = '1' then
              \state\ <= q_wait1637;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1635;
            end if;
          when pause_setII1657 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1653\ := \$arr1452_ptr_take\;
            if \$v1653\(0) = '1' then
              \state\ <= q_wait1652;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1650;
            end if;
          when pause_setII1668 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1665\ := \$arr1452_ptr_take\;
            if \$v1665\(0) = '1' then
              \state\ <= q_wait1664;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1662;
            end if;
          when pause_setII1704 =>
            \$arr1451_ptr_take\(0) := '0';
            \$208_y\ := \$224_x\;
            \$v1683\ := \$208_y\;
            \$v1684\ := \$v1683\(0 to 3);
            \$v1678\ := \$v1683\(4 to 35);
            case \$v1684\ is
            when "0001" =>
              \$26_a\ := \$v1678\(0 to 31);
              \$v1681\ := \$207_x\;
              \$v1682\ := \$v1681\(0 to 3);
              \$v1679\ := \$v1681\(4 to 35);
              case \$v1682\ is
              when "0001" =>
                b := \$v1679\(0 to 31);
                \$v1680\ := eclat_mult(\$26_a\ & b);
                \$209_result_after_f\ := "0001" & \$v1680\;
                \$v1677\ := \$arr1452_ptr_take\;
                if \$v1677\(0) = '1' then
                  \state\ <= q_wait1676;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1674;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("* arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811395\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("* arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811394\;
            end case;
          when pause_setII1772 =>
            \$arr1451_ptr_take\(0) := '0';
            \$207_x\ := \$270_x\;
            \$v1752\ := \$arr1452_ptr_take\;
            if \$v1752\(0) = '1' then
              \state\ <= q_wait1751;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1749;
            end if;
          when pause_setII1822 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v1820\ := \$arr1452_ptr_take\;
            if \$v1820\(0) = '1' then
              \state\ <= q_wait1819;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1817;
            end if;
          when pause_setII1839 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1835\ := \$arr1452_ptr_take\;
            if \$v1835\(0) = '1' then
              \state\ <= q_wait1834;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1832;
            end if;
          when pause_setII1850 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v1847\ := \$arr1452_ptr_take\;
            if \$v1847\(0) = '1' then
              \state\ <= q_wait1846;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1844;
            end if;
          when pause_setII1886 =>
            \$arr1451_ptr_take\(0) := '0';
            \$317_y\ := \$333_x\;
            \$v1865\ := \$317_y\;
            \$v1866\ := \$v1865\(0 to 3);
            \$v1860\ := \$v1865\(4 to 35);
            case \$v1866\ is
            when "0001" =>
              \$29_a\ := \$v1860\(0 to 31);
              \$v1863\ := \$316_x\;
              \$v1864\ := \$v1863\(0 to 3);
              \$v1861\ := \$v1863\(4 to 35);
              case \$v1864\ is
              when "0001" =>
                b := \$v1861\(0 to 31);
                \$v1862\ := eclat_sub(\$29_a\ & b);
                \$318_result_after_f\ := "0001" & \$v1862\;
                \$v1859\ := \$arr1452_ptr_take\;
                if \$v1859\(0) = '1' then
                  \state\ <= q_wait1858;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI1856;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("- arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811400\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("- arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811399\;
            end case;
          when pause_setII1954 =>
            \$arr1451_ptr_take\(0) := '0';
            \$316_x\ := \$379_x\;
            \$v1934\ := \$arr1452_ptr_take\;
            if \$v1934\(0) = '1' then
              \state\ <= q_wait1933;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1931;
            end if;
          when pause_setII2004 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2002\ := \$arr1452_ptr_take\;
            if \$v2002\(0) = '1' then
              \state\ <= q_wait2001;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1999;
            end if;
          when pause_setII2021 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2017\ := \$arr1452_ptr_take\;
            if \$v2017\(0) = '1' then
              \state\ <= q_wait2016;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2014;
            end if;
          when pause_setII2032 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2029\ := \$arr1452_ptr_take\;
            if \$v2029\(0) = '1' then
              \state\ <= q_wait2028;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2026;
            end if;
          when pause_setII2068 =>
            \$arr1451_ptr_take\(0) := '0';
            \$426_y\ := \$442_x\;
            \$v2047\ := \$426_y\;
            \$v2048\ := \$v2047\(0 to 3);
            \$v2042\ := \$v2047\(4 to 35);
            case \$v2048\ is
            when "0001" =>
              \$32_a\ := \$v2042\(0 to 31);
              \$v2045\ := \$425_x\;
              \$v2046\ := \$v2045\(0 to 3);
              \$v2043\ := \$v2045\(4 to 35);
              case \$v2046\ is
              when "0001" =>
                b := \$v2043\(0 to 31);
                \$v2044\ := eclat_add(\$32_a\ & b);
                \$427_result_after_f\ := "0001" & \$v2044\;
                \$v2041\ := \$arr1452_ptr_take\;
                if \$v2041\(0) = '1' then
                  \state\ <= q_wait2040;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2038;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("+ arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811405\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("+ arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811404\;
            end case;
          when pause_setII2136 =>
            \$arr1451_ptr_take\(0) := '0';
            \$425_x\ := \$488_x\;
            \$v2116\ := \$arr1452_ptr_take\;
            if \$v2116\(0) = '1' then
              \state\ <= q_wait2115;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2113;
            end if;
          when pause_setII2186 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2184\ := \$arr1452_ptr_take\;
            if \$v2184\(0) = '1' then
              \state\ <= q_wait2183;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2181;
            end if;
          when pause_setII2202 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2194\ := \$arr1452_ptr_take\;
            if \$v2194\(0) = '1' then
              \state\ <= q_wait2193;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2191;
            end if;
          when pause_setII2214 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2210\ := \$arr1452_ptr_take\;
            if \$v2210\(0) = '1' then
              \state\ <= q_wait2209;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2207;
            end if;
          when pause_setII2224 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2216\ := \$arr1451_ptr_take\;
            if \$v2216\(0) = '1' then
              \state\ <= q_wait2215;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2211\ := eclat_sub(\$82_i\ & "00000000000000000000000000000001");
              \$v2212\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2211\ & "0010" & \$82_i\ & "0001" & \$v2212\;
              \state\ <= pause_setI2213;
            end if;
          when pause_setII2259 =>
            \$arr1451_ptr_take\(0) := '0';
            \$53_y\ := \$540_x\;
            \$v2238\ := \$53_y\;
            \$v2239\ := \$v2238\(0 to 3);
            \$v2234\ := \$v2238\(4 to 35);
            case \$v2239\ is
            when "0001" =>
              \$35_a\ := \$v2234\(0 to 31);
              \$v2236\ := \$52_x\;
              \$v2237\ := \$v2236\(0 to 3);
              \$v2235\ := \$v2236\(4 to 35);
              case \$v2237\ is
              when "0001" =>
                b := \$v2235\(0 to 31);
                result := eclat_lt(\$35_a\ & b);
                \$v2233\ := \$arr1452_ptr_take\;
                if \$v2233\(0) = '1' then
                  \state\ <= q_wait2232;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2230;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("< arguments must be Ints"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$147_forever1811410\;
              end case;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("< arguments must be Ints"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811409\;
            end case;
          when pause_setII2327 =>
            \$arr1451_ptr_take\(0) := '0';
            \$52_x\ := \$586_x\;
            \$v2307\ := \$arr1452_ptr_take\;
            if \$v2307\(0) = '1' then
              \state\ <= q_wait2306;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2304;
            end if;
          when pause_setII2377 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2375\ := \$arr1452_ptr_take\;
            if \$v2375\(0) = '1' then
              \state\ <= q_wait2374;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2372;
            end if;
          when pause_setII2393 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2385\ := \$arr1452_ptr_take\;
            if \$v2385\(0) = '1' then
              \state\ <= q_wait2384;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2382;
            end if;
          when pause_setII2405 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2401\ := \$arr1452_ptr_take\;
            if \$v2401\(0) = '1' then
              \state\ <= q_wait2400;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2398;
            end if;
          when pause_setII2415 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2407\ := \$arr1451_ptr_take\;
            if \$v2407\(0) = '1' then
              \state\ <= q_wait2406;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2402\ := eclat_sub(\$635_i\ & "00000000000000000000000000000001");
              \$v2403\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2402\ & "0010" & \$635_i\ & "0001" & \$v2403\;
              \state\ <= pause_setI2404;
            end if;
          when pause_setII2453 =>
            \$arr1451_ptr_take\(0) := '0';
            \$633_y\ := \$642_x\;
            \$v2432\ := \$633_y\;
            \$v2433\ := \$v2432\(0 to 3);
            \$v2425\ := \$v2432\(4 to 35);
            case \$v2433\ is
            when "0010" =>
              ta := \$v2425\(0 to 31);
              \$v2427\ := \$632_x\;
              \$v2428\ := \$v2427\(0 to 3);
              \$v2426\ := \$v2427\(4 to 35);
              case \$v2428\ is
              when "0010" =>
                tb := \$v2426\(0 to 31);
                \$634_result\ := eclat_eq(ta & tb);
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              when others =>
                \$634_result\ := eclat_false;
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              end case;
            when "0001" =>
              ia := \$v2425\(0 to 31);
              \$v2430\ := \$632_x\;
              \$v2431\ := \$v2430\(0 to 3);
              \$v2429\ := \$v2430\(4 to 35);
              case \$v2431\ is
              when "0001" =>
                ib := \$v2429\(0 to 31);
                \$634_result\ := eclat_eq(ia & ib);
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              when others =>
                \$634_result\ := eclat_false;
                \$v2424\ := \$arr1452_ptr_take\;
                if \$v2424\(0) = '1' then
                  \state\ <= q_wait2423;
                else
                  \$arr1452_ptr_take\(0) := '1';
                  \$arr1452_ptr\ <= 1;
                  \state\ <= pause_getI2421;
                end if;
              end case;
            when others =>
              \$634_result\ := eclat_false;
              \$v2424\ := \$arr1452_ptr_take\;
              if \$v2424\(0) = '1' then
                \state\ <= q_wait2423;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI2421;
              end if;
            end case;
          when pause_setII2521 =>
            \$arr1451_ptr_take\(0) := '0';
            \$632_x\ := \$688_x\;
            \$v2501\ := \$arr1452_ptr_take\;
            if \$v2501\(0) = '1' then
              \state\ <= q_wait2500;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2498;
            end if;
          when pause_setII2571 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2569\ := \$arr1452_ptr_take\;
            if \$v2569\(0) = '1' then
              \state\ <= q_wait2568;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2566;
            end if;
          when pause_setII2581 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2579\ := \$arr1452_ptr_take\;
            if \$v2579\(0) = '1' then
              \state\ <= q_wait2578;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2576;
            end if;
          when pause_setII2593 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2589\ := \$arr1452_ptr_take\;
            if \$v2589\(0) = '1' then
              \state\ <= q_wait2588;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2586;
            end if;
          when pause_setII2597 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2595\ := \$arr1451_ptr_take\;
            if \$v2595\(0) = '1' then
              \state\ <= q_wait2594;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2590\ := eclat_sub(\$734_i\ & "00000000000000000000000000000001");
              \$v2591\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2590\ & "0010" & \$734_i\ & "0001" & \$v2591\;
              \state\ <= pause_setI2592;
            end if;
          when pause_setII2633 =>
            \$arr1451_ptr_take\(0) := '0';
            \$83_x\ := \$747_x\;
            \$v2612\ := \$83_x\;
            \$v2613\ := \$v2612\(0 to 3);
            \$v2607\ := \$v2612\(4 to 35);
            case \$v2613\ is
            when "0010" =>
              \$135_i\ := \$v2607\(0 to 31);
              \$v2611\ := \$arr1451_ptr_take\;
              if \$v2611\(0) = '1' then
                \state\ <= q_wait2610;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$135_i\));
                \state\ <= pause_getI2608;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811417\;
            end case;
          when pause_setII2701 =>
            \$arr1451_ptr_take\(0) := '0';
            \$55_x\ := \$793_x\;
            \$v2681\ := \$arr1452_ptr_take\;
            if \$v2681\(0) = '1' then
              \state\ <= q_wait2680;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2678;
            end if;
          when pause_setII2751 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2749\ := \$arr1452_ptr_take\;
            if \$v2749\(0) = '1' then
              \state\ <= q_wait2748;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2746;
            end if;
          when pause_setII2761 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2759\ := \$arr1452_ptr_take\;
            if \$v2759\(0) = '1' then
              \state\ <= q_wait2758;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2756;
            end if;
          when pause_setII2773 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2769\ := \$arr1452_ptr_take\;
            if \$v2769\(0) = '1' then
              \state\ <= q_wait2768;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2766;
            end if;
          when pause_setII2777 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2775\ := \$arr1451_ptr_take\;
            if \$v2775\(0) = '1' then
              \state\ <= q_wait2774;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2770\ := eclat_sub(\$841_i\ & "00000000000000000000000000000001");
              \$v2771\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2770\ & "0010" & \$841_i\ & "0001" & \$v2771\;
              \state\ <= pause_setI2772;
            end if;
          when pause_setII2813 =>
            \$arr1451_ptr_take\(0) := '0';
            \$851_x\ := \$856_x\;
            \$v2792\ := \$851_x\;
            \$v2793\ := \$v2792\(0 to 3);
            \$v2787\ := \$v2792\(4 to 35);
            case \$v2793\ is
            when "0010" =>
              \$852_i\ := \$v2787\(0 to 31);
              \$v2791\ := \$arr1451_ptr_take\;
              if \$v2791\(0) = '1' then
                \state\ <= q_wait2790;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$852_i\));
                \state\ <= pause_getI2788;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811421\;
            end case;
          when pause_setII2881 =>
            \$arr1451_ptr_take\(0) := '0';
            \$839_x\ := \$902_x\;
            \$v2861\ := \$arr1452_ptr_take\;
            if \$v2861\(0) = '1' then
              \state\ <= q_wait2860;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2858;
            end if;
          when pause_setII2931 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v2929\ := \$arr1452_ptr_take\;
            if \$v2929\(0) = '1' then
              \state\ <= q_wait2928;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2926;
            end if;
          when pause_setII2941 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2939\ := \$arr1452_ptr_take\;
            if \$v2939\(0) = '1' then
              \state\ <= q_wait2938;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2936;
            end if;
          when pause_setII2953 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2949\ := \$arr1452_ptr_take\;
            if \$v2949\(0) = '1' then
              \state\ <= q_wait2948;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2946;
            end if;
          when pause_setII2957 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v2955\ := \$arr1451_ptr_take\;
            if \$v2955\(0) = '1' then
              \state\ <= q_wait2954;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2950\ := eclat_sub(\$950_i\ & "00000000000000000000000000000001");
              \$v2951\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2950\ & "0010" & \$950_i\ & "0001" & \$v2951\;
              \state\ <= pause_setI2952;
            end if;
          when pause_setII2993 =>
            \$arr1451_ptr_take\(0) := '0';
            \$960_x\ := \$965_x\;
            \$v2972\ := \$960_x\;
            \$v2973\ := \$v2972\(0 to 3);
            \$v2967\ := \$v2972\(4 to 35);
            case \$v2973\ is
            when "0010" =>
              \$961_i\ := \$v2967\(0 to 31);
              \$v2971\ := \$arr1451_ptr_take\;
              if \$v2971\(0) = '1' then
                \state\ <= q_wait2970;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$961_i\));
                \state\ <= pause_getI2968;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811425\;
            end case;
          when pause_setII3061 =>
            \$arr1451_ptr_take\(0) := '0';
            \$948_x\ := \$1011_x\;
            \$v3041\ := \$arr1452_ptr_take\;
            if \$v3041\(0) = '1' then
              \state\ <= q_wait3040;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3038;
            end if;
          when pause_setII3111 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3109\ := \$arr1452_ptr_take\;
            if \$v3109\(0) = '1' then
              \state\ <= q_wait3108;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3106;
            end if;
          when pause_setII3128 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3124\ := \$arr1452_ptr_take\;
            if \$v3124\(0) = '1' then
              \state\ <= q_wait3123;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3121;
            end if;
          when pause_setII3139 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3136\ := \$arr1452_ptr_take\;
            if \$v3136\(0) = '1' then
              \state\ <= q_wait3135;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3133;
            end if;
          when pause_setII3175 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1074_x\ := \$1079_x\;
            \$v3154\ := \$1074_x\;
            \$v3155\ := \$v3154\(0 to 3);
            \$v3149\ := \$v3154\(4 to 35);
            case \$v3155\ is
            when "0010" =>
              \$1075_i\ := \$v3149\(0 to 31);
              \$v3153\ := \$arr1451_ptr_take\;
              if \$v3153\(0) = '1' then
                \state\ <= q_wait3152;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1075_i\));
                \state\ <= pause_getI3150;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811429\;
            end case;
          when pause_setII3225 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3223\ := \$arr1452_ptr_take\;
            if \$v3223\(0) = '1' then
              \state\ <= q_wait3222;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3220;
            end if;
          when pause_setII3242 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3238\ := \$arr1452_ptr_take\;
            if \$v3238\(0) = '1' then
              \state\ <= q_wait3237;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3235;
            end if;
          when pause_setII3253 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3250\ := \$arr1452_ptr_take\;
            if \$v3250\(0) = '1' then
              \state\ <= q_wait3249;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3247;
            end if;
          when pause_setII3289 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1143_x\ := \$1148_x\;
            \$v3268\ := \$1143_x\;
            \$v3269\ := \$v3268\(0 to 3);
            \$v3263\ := \$v3268\(4 to 35);
            case \$v3269\ is
            when "0010" =>
              \$1144_i\ := \$v3263\(0 to 31);
              \$v3267\ := \$arr1451_ptr_take\;
              if \$v3267\(0) = '1' then
                \state\ <= q_wait3266;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1144_i\));
                \state\ <= pause_getI3264;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811432\;
            end case;
          when pause_setII3339 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3337\ := \$arr1452_ptr_take\;
            if \$v3337\(0) = '1' then
              \state\ <= q_wait3336;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3334;
            end if;
          when pause_setII3356 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3352\ := \$arr1452_ptr_take\;
            if \$v3352\(0) = '1' then
              \state\ <= q_wait3351;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3349;
            end if;
          when pause_setII3367 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3364\ := \$arr1452_ptr_take\;
            if \$v3364\(0) = '1' then
              \state\ <= q_wait3363;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3361;
            end if;
          when pause_setII3403 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1212_x\ := \$1217_x\;
            \$v3382\ := \$1212_x\;
            \$v3383\ := \$v3382\(0 to 3);
            \$v3377\ := \$v3382\(4 to 35);
            case \$v3383\ is
            when "0010" =>
              \$1213_i\ := \$v3377\(0 to 31);
              \$v3381\ := \$arr1451_ptr_take\;
              if \$v3381\(0) = '1' then
                \state\ <= q_wait3380;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1213_i\));
                \state\ <= pause_getI3378;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811435\;
            end case;
          when pause_setII3453 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3451\ := \$arr1452_ptr_take\;
            if \$v3451\(0) = '1' then
              \state\ <= q_wait3450;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3448;
            end if;
          when pause_setII3463 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3461\ := \$arr1452_ptr_take\;
            if \$v3461\(0) = '1' then
              \state\ <= q_wait3460;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3458;
            end if;
          when pause_setII3475 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3471\ := \$arr1452_ptr_take\;
            if \$v3471\(0) = '1' then
              \state\ <= q_wait3470;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3468;
            end if;
          when pause_setII3479 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3477\ := \$arr1451_ptr_take\;
            if \$v3477\(0) = '1' then
              \state\ <= q_wait3476;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3472\ := eclat_sub(\$1263_i\ & "00000000000000000000000000000001");
              \$v3473\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3472\ & "0010" & \$1263_i\ & "0001" & \$v3473\;
              \state\ <= pause_setI3474;
            end if;
          when pause_setII3517 =>
            \$arr1451_ptr_take\(0) := '0';
            \$73_result\ := \$1270_x\;
            \$v3496\ := \$73_result\;
            \$v3497\ := \$v3496\(0 to 3);
            \$v3489\ := \$v3496\(4 to 35);
            case \$v3497\ is
            when "0010" =>
              \$v3490\ := "00000000000000000000000000000000";
              \$v3491\ := "00000000000000000000000000000000";
              \$v3492\ := "00000000000000000000000000000101";
              \$74_result_after_f\ := "0001" & \$v3490\ & "0001" & \$v3491\ & "0001" & \$v3492\;
              \$v3488\ := \$arr1452_ptr_take\;
              if \$v3488\(0) = '1' then
                \state\ <= q_wait3487;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3485;
              end if;
            when others =>
              \$v3493\ := "00000000000000000000000000000001";
              \$v3494\ := "00000000000000000000000000000010";
              \$v3495\ := "00000000000000000000000000000101";
              \$74_result_after_f\ := "0010" & \$v3493\ & "0010" & \$v3494\ & "0001" & \$v3495\;
              \$v3488\ := \$arr1452_ptr_take\;
              if \$v3488\(0) = '1' then
                \state\ <= q_wait3487;
              else
                \$arr1452_ptr_take\(0) := '1';
                \$arr1452_ptr\ <= 1;
                \state\ <= pause_getI3485;
              end if;
            end case;
          when pause_setII3567 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3565\ := \$arr1452_ptr_take\;
            if \$v3565\(0) = '1' then
              \state\ <= q_wait3564;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3562;
            end if;
          when pause_setII3578 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3575\ := \$arr1452_ptr_take\;
            if \$v3575\(0) = '1' then
              \state\ <= q_wait3574;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3572;
            end if;
          when pause_setII3590 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3586\ := \$arr1452_ptr_take\;
            if \$v3586\(0) = '1' then
              \state\ <= q_wait3585;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3583;
            end if;
          when pause_setII3595 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3592\ := \$arr1451_ptr_take\;
            if \$v3592\(0) = '1' then
              \state\ <= q_wait3591;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3587\ := eclat_sub(\$1316_i\ & "00000000000000000000000000000001");
              \$v3588\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3587\ & "0010" & \$1316_i\ & "0001" & \$v3588\;
              \state\ <= pause_setI3589;
            end if;
          when pause_setII3640 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1332_x\ := \$1337_x\;
            \$v3619\ := \$1332_x\;
            \$v3620\ := \$v3619\(0 to 3);
            \$v3614\ := \$v3619\(4 to 35);
            case \$v3620\ is
            when "0010" =>
              \$1333_i\ := \$v3614\(0 to 31);
              \$v3618\ := \$arr1451_ptr_take\;
              if \$v3618\(0) = '1' then
                \state\ <= q_wait3617;
              else
                \$arr1451_ptr_take\(0) := '1';
                \$arr1451_ptr\ <= to_integer(unsigned(\$1333_i\));
                \state\ <= pause_getI3615;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_rib expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$147_forever1811440\;
            end case;
          when pause_setII3690 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3688\ := \$arr1452_ptr_take\;
            if \$v3688\(0) = '1' then
              \state\ <= q_wait3687;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3685;
            end if;
          when pause_setII3707 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3703\ := \$arr1452_ptr_take\;
            if \$v3703\(0) = '1' then
              \state\ <= q_wait3702;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3700;
            end if;
          when pause_setII3718 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3715\ := \$arr1452_ptr_take\;
            if \$v3715\(0) = '1' then
              \state\ <= q_wait3714;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3712;
            end if;
          when pause_setII3747 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3727\ := \$arr1452_ptr_take\;
            if \$v3727\(0) = '1' then
              \state\ <= q_wait3726;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3724;
            end if;
          when pause_setII3815 =>
            \$arr1451_ptr_take\(0) := '0';
            \$1383_x\ := \$1442_x\;
            \$v3795\ := \$arr1452_ptr_take\;
            if \$v3795\(0) = '1' then
              \state\ <= q_wait3794;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3792;
            end if;
          when pause_setII3865 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3863\ := \$arr1452_ptr_take\;
            if \$v3863\(0) = '1' then
              \state\ <= q_wait3862;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3860;
            end if;
          when pause_setII3882 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3878\ := \$arr1452_ptr_take\;
            if \$v3878\(0) = '1' then
              \state\ <= q_wait3877;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3875;
            end if;
          when pause_setII3893 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3890\ := \$arr1452_ptr_take\;
            if \$v3890\(0) = '1' then
              \state\ <= q_wait3889;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3887;
            end if;
          when pause_setII3922 =>
            \$arr1451_ptr_take\(0) := '0';
            \$76_result\ := \$1499_x\;
            \$v3902\ := \$arr1452_ptr_take\;
            if \$v3902\(0) = '1' then
              \state\ <= q_wait3901;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3899;
            end if;
          when pause_setII3972 =>
            \$arr1453_ptr_take\(0) := '0';
            \$v3970\ := \$arr1452_ptr_take\;
            if \$v3970\(0) = '1' then
              \state\ <= q_wait3969;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3967;
            end if;
          when pause_setII3982 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3980\ := \$arr1452_ptr_take\;
            if \$v3980\(0) = '1' then
              \state\ <= q_wait3979;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3977;
            end if;
          when pause_setII3994 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3990\ := \$arr1452_ptr_take\;
            if \$v3990\(0) = '1' then
              \state\ <= q_wait3989;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3987;
            end if;
          when pause_setII3998 =>
            \$arr1451_ptr_take\(0) := '0';
            \$v3996\ := \$arr1451_ptr_take\;
            if \$v3996\(0) = '1' then
              \state\ <= q_wait3995;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3991\ := eclat_sub(\$1545_i\ & "00000000000000000000000000000001");
              \$v3992\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3991\ & "0010" & \$1545_i\ & "0001" & \$v3992\;
              \state\ <= pause_setI3993;
            end if;
          when pause_setII4027 =>
            \$arr1451_ptr_take\(0) := '0';
            \$67_z\ := \$1552_x\;
            \$v4007\ := \$arr1452_ptr_take\;
            if \$v4007\(0) = '1' then
              \state\ <= q_wait4006;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4004;
            end if;
          when pause_setII4095 =>
            \$arr1451_ptr_take\(0) := '0';
            \$66_y\ := \$1598_x\;
            \$v4075\ := \$arr1452_ptr_take\;
            if \$v4075\(0) = '1' then
              \state\ <= q_wait4074;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4072;
            end if;
          when pause_setII4163 =>
            \$arr1451_ptr_take\(0) := '0';
            \$65_x\ := \$1644_x\;
            \$v4143\ := \$arr1452_ptr_take\;
            if \$v4143\(0) = '1' then
              \state\ <= q_wait4142;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4140;
            end if;
          when pause_setII4222 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4220\ := \$arr1452_ptr_take\;
            if \$v4220\(0) = '1' then
              \state\ <= q_wait4219;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4217;
            end if;
          when pause_setII4226 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4224\ := \$arr1452_ptr_take\;
            if \$v4224\(0) = '1' then
              \state\ <= q_wait4223;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 4;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= pos;
              \state\ <= pause_setI4221;
            end if;
          when pause_setII4230 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4228\ := \$arr1452_ptr_take\;
            if \$v4228\(0) = '1' then
              \state\ <= q_wait4227;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 3;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= stbl;
              \state\ <= pause_setI4225;
            end if;
          when pause_setII4234 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4232\ := \$arr1452_ptr_take\;
            if \$v4232\(0) = '1' then
              \state\ <= q_wait4231;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 2;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= st;
              \state\ <= pause_setI4229;
            end if;
          when pause_setII4238 =>
            \$arr1452_ptr_take\(0) := '0';
            \$v4236\ := \$arr1452_ptr_take\;
            if \$v4236\(0) = '1' then
              \state\ <= q_wait4235;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 1;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= sp;
              \state\ <= pause_setI4233;
            end if;
          when q_wait1459 =>
            \$v1460\ := \$arr1453_ptr_take\;
            if \$v1460\(0) = '1' then
              \state\ <= q_wait1459;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 17;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v120\;
              \state\ <= pause_setI1457;
            end if;
          when q_wait1466 =>
            \$v1467\ := \$arr1452_ptr_take\;
            if \$v1467\(0) = '1' then
              \state\ <= q_wait1466;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1464;
            end if;
          when q_wait1470 =>
            \$v1471\ := \$arr1452_ptr_take\;
            if \$v1471\(0) = '1' then
              \state\ <= q_wait1470;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1468;
            end if;
          when q_wait1476 =>
            \$v1477\ := \$arr1451_ptr_take\;
            if \$v1477\(0) = '1' then
              \state\ <= q_wait1476;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1472\ := "00000000000000000000000000000000";
              \$v1473\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$71_result_after_f\ & "0001" & \$v1472\ & "0001" & \$v1473\;
              \state\ <= pause_setI1474;
            end if;
          when q_wait1482 =>
            \$v1483\ := \$arr1452_ptr_take\;
            if \$v1483\(0) = '1' then
              \state\ <= q_wait1482;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1480;
            end if;
          when q_wait1487 =>
            \$v1488\ := \$arr1451_ptr_take\;
            if \$v1488\(0) = '1' then
              \state\ <= q_wait1487;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1484\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$81_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$71_result_after_f\ & "0010" & \$81_i\ & "0001" & \$v1484\;
              \state\ <= pause_setI1485;
            end if;
          when q_wait1494 =>
            \$v1495\ := \$arr1452_ptr_take\;
            if \$v1495\(0) = '1' then
              \state\ <= q_wait1494;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1492;
            end if;
          when q_wait1510 =>
            \$v1511\ := \$arr1451_ptr_take\;
            if \$v1511\(0) = '1' then
              \state\ <= q_wait1510;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v40\));
              \state\ <= pause_getI1508;
            end if;
          when q_wait1515 =>
            \$v1516\ := \$arr1452_ptr_take\;
            if \$v1516\(0) = '1' then
              \state\ <= q_wait1515;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1513;
            end if;
          when q_wait1519 =>
            \$v1520\ := \$arr1452_ptr_take\;
            if \$v1520\(0) = '1' then
              \state\ <= q_wait1519;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1517;
            end if;
          when q_wait1523 =>
            \$v1524\ := \$arr1451_ptr_take\;
            if \$v1524\(0) = '1' then
              \state\ <= q_wait1523;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$v37\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$v38\;
              \state\ <= pause_setI1521;
            end if;
          when q_wait1528 =>
            \$v1529\ := \$arr1451_ptr_take\;
            if \$v1529\(0) = '1' then
              \state\ <= q_wait1528;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v32\));
              \state\ <= pause_getI1526;
            end if;
          when q_wait1533 =>
            \$v1534\ := \$arr1452_ptr_take\;
            if \$v1534\(0) = '1' then
              \state\ <= q_wait1533;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1531;
            end if;
          when q_wait1537 =>
            \$v1538\ := \$arr1451_ptr_take\;
            if \$v1538\(0) = '1' then
              \state\ <= q_wait1537;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v29\));
              \state\ <= pause_getI1535;
            end if;
          when q_wait1542 =>
            \$v1543\ := \$arr1452_ptr_take\;
            if \$v1543\(0) = '1' then
              \state\ <= q_wait1542;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1540;
            end if;
          when q_wait1547 =>
            \$v1548\ := \$arr1452_ptr_take\;
            if \$v1548\(0) = '1' then
              \state\ <= q_wait1547;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1545;
            end if;
          when q_wait1555 =>
            \$v1556\ := \$arr1451_ptr_take\;
            if \$v1556\(0) = '1' then
              \state\ <= q_wait1555;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v23\));
              \state\ <= pause_getI1553;
            end if;
          when q_wait1560 =>
            \$v1561\ := \$arr1452_ptr_take\;
            if \$v1561\(0) = '1' then
              \state\ <= q_wait1560;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1558;
            end if;
          when q_wait1564 =>
            \$v1565\ := \$arr1451_ptr_take\;
            if \$v1565\(0) = '1' then
              \state\ <= q_wait1564;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v20\));
              \state\ <= pause_getI1562;
            end if;
          when q_wait1569 =>
            \$v1570\ := \$arr1452_ptr_take\;
            if \$v1570\(0) = '1' then
              \state\ <= q_wait1569;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1567;
            end if;
          when q_wait1578 =>
            \$v1579\ := \$arr1451_ptr_take\;
            if \$v1579\(0) = '1' then
              \state\ <= q_wait1578;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$191\));
              \state\ <= pause_getI1576;
            end if;
          when q_wait1583 =>
            \$v1584\ := \$arr1452_ptr_take\;
            if \$v1584\(0) = '1' then
              \state\ <= q_wait1583;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1581;
            end if;
          when q_wait1587 =>
            \$v1588\ := \$arr1452_ptr_take\;
            if \$v1588\(0) = '1' then
              \state\ <= q_wait1587;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1585;
            end if;
          when q_wait1591 =>
            \$v1592\ := \$arr1451_ptr_take\;
            if \$v1592\(0) = '1' then
              \state\ <= q_wait1591;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$163\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$164\;
              \state\ <= pause_setI1589;
            end if;
          when q_wait1596 =>
            \$v1597\ := \$arr1451_ptr_take\;
            if \$v1597\(0) = '1' then
              \state\ <= q_wait1596;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$171\));
              \state\ <= pause_getI1594;
            end if;
          when q_wait1601 =>
            \$v1602\ := \$arr1452_ptr_take\;
            if \$v1602\(0) = '1' then
              \state\ <= q_wait1601;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1599;
            end if;
          when q_wait1605 =>
            \$v1606\ := \$arr1451_ptr_take\;
            if \$v1606\(0) = '1' then
              \state\ <= q_wait1605;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$177\));
              \state\ <= pause_getI1603;
            end if;
          when q_wait1610 =>
            \$v1611\ := \$arr1452_ptr_take\;
            if \$v1611\(0) = '1' then
              \state\ <= q_wait1610;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1608;
            end if;
          when q_wait1615 =>
            \$v1616\ := \$arr1452_ptr_take\;
            if \$v1616\(0) = '1' then
              \state\ <= q_wait1615;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1613;
            end if;
          when q_wait1623 =>
            \$v1624\ := \$arr1451_ptr_take\;
            if \$v1624\(0) = '1' then
              \state\ <= q_wait1623;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$199\));
              \state\ <= pause_getI1621;
            end if;
          when q_wait1628 =>
            \$v1629\ := \$arr1452_ptr_take\;
            if \$v1629\(0) = '1' then
              \state\ <= q_wait1628;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1626;
            end if;
          when q_wait1632 =>
            \$v1633\ := \$arr1451_ptr_take\;
            if \$v1633\(0) = '1' then
              \state\ <= q_wait1632;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$205\));
              \state\ <= pause_getI1630;
            end if;
          when q_wait1637 =>
            \$v1638\ := \$arr1452_ptr_take\;
            if \$v1638\(0) = '1' then
              \state\ <= q_wait1637;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1635;
            end if;
          when q_wait1641 =>
            \$v1642\ := \$arr1453_ptr_take\;
            if \$v1642\(0) = '1' then
              \state\ <= q_wait1641;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 16;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v117\;
              \state\ <= pause_setI1639;
            end if;
          when q_wait1648 =>
            \$v1649\ := \$arr1452_ptr_take\;
            if \$v1649\(0) = '1' then
              \state\ <= q_wait1648;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1646;
            end if;
          when q_wait1652 =>
            \$v1653\ := \$arr1452_ptr_take\;
            if \$v1653\(0) = '1' then
              \state\ <= q_wait1652;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1650;
            end if;
          when q_wait1658 =>
            \$v1659\ := \$arr1451_ptr_take\;
            if \$v1659\(0) = '1' then
              \state\ <= q_wait1658;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1654\ := "00000000000000000000000000000000";
              \$v1655\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$209_result_after_f\ & "0001" & \$v1654\ & "0001" & \$v1655\;
              \state\ <= pause_setI1656;
            end if;
          when q_wait1664 =>
            \$v1665\ := \$arr1452_ptr_take\;
            if \$v1665\(0) = '1' then
              \state\ <= q_wait1664;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1662;
            end if;
          when q_wait1669 =>
            \$v1670\ := \$arr1451_ptr_take\;
            if \$v1670\(0) = '1' then
              \state\ <= q_wait1669;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1666\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$210_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$209_result_after_f\ & "0010" & \$210_i\ & "0001" & \$v1666\;
              \state\ <= pause_setI1667;
            end if;
          when q_wait1676 =>
            \$v1677\ := \$arr1452_ptr_take\;
            if \$v1677\(0) = '1' then
              \state\ <= q_wait1676;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1674;
            end if;
          when q_wait1692 =>
            \$v1693\ := \$arr1451_ptr_take\;
            if \$v1693\(0) = '1' then
              \state\ <= q_wait1692;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$254\));
              \state\ <= pause_getI1690;
            end if;
          when q_wait1697 =>
            \$v1698\ := \$arr1452_ptr_take\;
            if \$v1698\(0) = '1' then
              \state\ <= q_wait1697;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1695;
            end if;
          when q_wait1701 =>
            \$v1702\ := \$arr1452_ptr_take\;
            if \$v1702\(0) = '1' then
              \state\ <= q_wait1701;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1699;
            end if;
          when q_wait1705 =>
            \$v1706\ := \$arr1451_ptr_take\;
            if \$v1706\(0) = '1' then
              \state\ <= q_wait1705;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$226\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$227\;
              \state\ <= pause_setI1703;
            end if;
          when q_wait1710 =>
            \$v1711\ := \$arr1451_ptr_take\;
            if \$v1711\(0) = '1' then
              \state\ <= q_wait1710;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$234\));
              \state\ <= pause_getI1708;
            end if;
          when q_wait1715 =>
            \$v1716\ := \$arr1452_ptr_take\;
            if \$v1716\(0) = '1' then
              \state\ <= q_wait1715;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1713;
            end if;
          when q_wait1719 =>
            \$v1720\ := \$arr1451_ptr_take\;
            if \$v1720\(0) = '1' then
              \state\ <= q_wait1719;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$240\));
              \state\ <= pause_getI1717;
            end if;
          when q_wait1724 =>
            \$v1725\ := \$arr1452_ptr_take\;
            if \$v1725\(0) = '1' then
              \state\ <= q_wait1724;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1722;
            end if;
          when q_wait1729 =>
            \$v1730\ := \$arr1452_ptr_take\;
            if \$v1730\(0) = '1' then
              \state\ <= q_wait1729;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1727;
            end if;
          when q_wait1737 =>
            \$v1738\ := \$arr1451_ptr_take\;
            if \$v1738\(0) = '1' then
              \state\ <= q_wait1737;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$262\));
              \state\ <= pause_getI1735;
            end if;
          when q_wait1742 =>
            \$v1743\ := \$arr1452_ptr_take\;
            if \$v1743\(0) = '1' then
              \state\ <= q_wait1742;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1740;
            end if;
          when q_wait1746 =>
            \$v1747\ := \$arr1451_ptr_take\;
            if \$v1747\(0) = '1' then
              \state\ <= q_wait1746;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$268\));
              \state\ <= pause_getI1744;
            end if;
          when q_wait1751 =>
            \$v1752\ := \$arr1452_ptr_take\;
            if \$v1752\(0) = '1' then
              \state\ <= q_wait1751;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1749;
            end if;
          when q_wait1760 =>
            \$v1761\ := \$arr1451_ptr_take\;
            if \$v1761\(0) = '1' then
              \state\ <= q_wait1760;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$300\));
              \state\ <= pause_getI1758;
            end if;
          when q_wait1765 =>
            \$v1766\ := \$arr1452_ptr_take\;
            if \$v1766\(0) = '1' then
              \state\ <= q_wait1765;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1763;
            end if;
          when q_wait1769 =>
            \$v1770\ := \$arr1452_ptr_take\;
            if \$v1770\(0) = '1' then
              \state\ <= q_wait1769;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1767;
            end if;
          when q_wait1773 =>
            \$v1774\ := \$arr1451_ptr_take\;
            if \$v1774\(0) = '1' then
              \state\ <= q_wait1773;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$272\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$273\;
              \state\ <= pause_setI1771;
            end if;
          when q_wait1778 =>
            \$v1779\ := \$arr1451_ptr_take\;
            if \$v1779\(0) = '1' then
              \state\ <= q_wait1778;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$280\));
              \state\ <= pause_getI1776;
            end if;
          when q_wait1783 =>
            \$v1784\ := \$arr1452_ptr_take\;
            if \$v1784\(0) = '1' then
              \state\ <= q_wait1783;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1781;
            end if;
          when q_wait1787 =>
            \$v1788\ := \$arr1451_ptr_take\;
            if \$v1788\(0) = '1' then
              \state\ <= q_wait1787;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$286\));
              \state\ <= pause_getI1785;
            end if;
          when q_wait1792 =>
            \$v1793\ := \$arr1452_ptr_take\;
            if \$v1793\(0) = '1' then
              \state\ <= q_wait1792;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1790;
            end if;
          when q_wait1797 =>
            \$v1798\ := \$arr1452_ptr_take\;
            if \$v1798\(0) = '1' then
              \state\ <= q_wait1797;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1795;
            end if;
          when q_wait1805 =>
            \$v1806\ := \$arr1451_ptr_take\;
            if \$v1806\(0) = '1' then
              \state\ <= q_wait1805;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$308\));
              \state\ <= pause_getI1803;
            end if;
          when q_wait1810 =>
            \$v1811\ := \$arr1452_ptr_take\;
            if \$v1811\(0) = '1' then
              \state\ <= q_wait1810;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1808;
            end if;
          when q_wait1814 =>
            \$v1815\ := \$arr1451_ptr_take\;
            if \$v1815\(0) = '1' then
              \state\ <= q_wait1814;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$314\));
              \state\ <= pause_getI1812;
            end if;
          when q_wait1819 =>
            \$v1820\ := \$arr1452_ptr_take\;
            if \$v1820\(0) = '1' then
              \state\ <= q_wait1819;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1817;
            end if;
          when q_wait1823 =>
            \$v1824\ := \$arr1453_ptr_take\;
            if \$v1824\(0) = '1' then
              \state\ <= q_wait1823;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 15;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v114\;
              \state\ <= pause_setI1821;
            end if;
          when q_wait1830 =>
            \$v1831\ := \$arr1452_ptr_take\;
            if \$v1831\(0) = '1' then
              \state\ <= q_wait1830;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1828;
            end if;
          when q_wait1834 =>
            \$v1835\ := \$arr1452_ptr_take\;
            if \$v1835\(0) = '1' then
              \state\ <= q_wait1834;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1832;
            end if;
          when q_wait1840 =>
            \$v1841\ := \$arr1451_ptr_take\;
            if \$v1841\(0) = '1' then
              \state\ <= q_wait1840;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1836\ := "00000000000000000000000000000000";
              \$v1837\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$318_result_after_f\ & "0001" & \$v1836\ & "0001" & \$v1837\;
              \state\ <= pause_setI1838;
            end if;
          when q_wait1846 =>
            \$v1847\ := \$arr1452_ptr_take\;
            if \$v1847\(0) = '1' then
              \state\ <= q_wait1846;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1844;
            end if;
          when q_wait1851 =>
            \$v1852\ := \$arr1451_ptr_take\;
            if \$v1852\(0) = '1' then
              \state\ <= q_wait1851;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v1848\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$319_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$318_result_after_f\ & "0010" & \$319_i\ & "0001" & \$v1848\;
              \state\ <= pause_setI1849;
            end if;
          when q_wait1858 =>
            \$v1859\ := \$arr1452_ptr_take\;
            if \$v1859\(0) = '1' then
              \state\ <= q_wait1858;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1856;
            end if;
          when q_wait1874 =>
            \$v1875\ := \$arr1451_ptr_take\;
            if \$v1875\(0) = '1' then
              \state\ <= q_wait1874;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$363\));
              \state\ <= pause_getI1872;
            end if;
          when q_wait1879 =>
            \$v1880\ := \$arr1452_ptr_take\;
            if \$v1880\(0) = '1' then
              \state\ <= q_wait1879;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1877;
            end if;
          when q_wait1883 =>
            \$v1884\ := \$arr1452_ptr_take\;
            if \$v1884\(0) = '1' then
              \state\ <= q_wait1883;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1881;
            end if;
          when q_wait1887 =>
            \$v1888\ := \$arr1451_ptr_take\;
            if \$v1888\(0) = '1' then
              \state\ <= q_wait1887;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$335\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$336\;
              \state\ <= pause_setI1885;
            end if;
          when q_wait1892 =>
            \$v1893\ := \$arr1451_ptr_take\;
            if \$v1893\(0) = '1' then
              \state\ <= q_wait1892;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$343\));
              \state\ <= pause_getI1890;
            end if;
          when q_wait1897 =>
            \$v1898\ := \$arr1452_ptr_take\;
            if \$v1898\(0) = '1' then
              \state\ <= q_wait1897;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1895;
            end if;
          when q_wait1901 =>
            \$v1902\ := \$arr1451_ptr_take\;
            if \$v1902\(0) = '1' then
              \state\ <= q_wait1901;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$349\));
              \state\ <= pause_getI1899;
            end if;
          when q_wait1906 =>
            \$v1907\ := \$arr1452_ptr_take\;
            if \$v1907\(0) = '1' then
              \state\ <= q_wait1906;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1904;
            end if;
          when q_wait1911 =>
            \$v1912\ := \$arr1452_ptr_take\;
            if \$v1912\(0) = '1' then
              \state\ <= q_wait1911;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1909;
            end if;
          when q_wait1919 =>
            \$v1920\ := \$arr1451_ptr_take\;
            if \$v1920\(0) = '1' then
              \state\ <= q_wait1919;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$371\));
              \state\ <= pause_getI1917;
            end if;
          when q_wait1924 =>
            \$v1925\ := \$arr1452_ptr_take\;
            if \$v1925\(0) = '1' then
              \state\ <= q_wait1924;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1922;
            end if;
          when q_wait1928 =>
            \$v1929\ := \$arr1451_ptr_take\;
            if \$v1929\(0) = '1' then
              \state\ <= q_wait1928;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$377\));
              \state\ <= pause_getI1926;
            end if;
          when q_wait1933 =>
            \$v1934\ := \$arr1452_ptr_take\;
            if \$v1934\(0) = '1' then
              \state\ <= q_wait1933;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1931;
            end if;
          when q_wait1942 =>
            \$v1943\ := \$arr1451_ptr_take\;
            if \$v1943\(0) = '1' then
              \state\ <= q_wait1942;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$409\));
              \state\ <= pause_getI1940;
            end if;
          when q_wait1947 =>
            \$v1948\ := \$arr1452_ptr_take\;
            if \$v1948\(0) = '1' then
              \state\ <= q_wait1947;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1945;
            end if;
          when q_wait1951 =>
            \$v1952\ := \$arr1452_ptr_take\;
            if \$v1952\(0) = '1' then
              \state\ <= q_wait1951;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1949;
            end if;
          when q_wait1955 =>
            \$v1956\ := \$arr1451_ptr_take\;
            if \$v1956\(0) = '1' then
              \state\ <= q_wait1955;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$381\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$382\;
              \state\ <= pause_setI1953;
            end if;
          when q_wait1960 =>
            \$v1961\ := \$arr1451_ptr_take\;
            if \$v1961\(0) = '1' then
              \state\ <= q_wait1960;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$389\));
              \state\ <= pause_getI1958;
            end if;
          when q_wait1965 =>
            \$v1966\ := \$arr1452_ptr_take\;
            if \$v1966\(0) = '1' then
              \state\ <= q_wait1965;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1963;
            end if;
          when q_wait1969 =>
            \$v1970\ := \$arr1451_ptr_take\;
            if \$v1970\(0) = '1' then
              \state\ <= q_wait1969;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$395\));
              \state\ <= pause_getI1967;
            end if;
          when q_wait1974 =>
            \$v1975\ := \$arr1452_ptr_take\;
            if \$v1975\(0) = '1' then
              \state\ <= q_wait1974;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1972;
            end if;
          when q_wait1979 =>
            \$v1980\ := \$arr1452_ptr_take\;
            if \$v1980\(0) = '1' then
              \state\ <= q_wait1979;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1977;
            end if;
          when q_wait1987 =>
            \$v1988\ := \$arr1451_ptr_take\;
            if \$v1988\(0) = '1' then
              \state\ <= q_wait1987;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$417\));
              \state\ <= pause_getI1985;
            end if;
          when q_wait1992 =>
            \$v1993\ := \$arr1452_ptr_take\;
            if \$v1993\(0) = '1' then
              \state\ <= q_wait1992;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1990;
            end if;
          when q_wait1996 =>
            \$v1997\ := \$arr1451_ptr_take\;
            if \$v1997\(0) = '1' then
              \state\ <= q_wait1996;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$423\));
              \state\ <= pause_getI1994;
            end if;
          when q_wait2001 =>
            \$v2002\ := \$arr1452_ptr_take\;
            if \$v2002\(0) = '1' then
              \state\ <= q_wait2001;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI1999;
            end if;
          when q_wait2005 =>
            \$v2006\ := \$arr1453_ptr_take\;
            if \$v2006\(0) = '1' then
              \state\ <= q_wait2005;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 14;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v111\;
              \state\ <= pause_setI2003;
            end if;
          when q_wait2012 =>
            \$v2013\ := \$arr1452_ptr_take\;
            if \$v2013\(0) = '1' then
              \state\ <= q_wait2012;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2010;
            end if;
          when q_wait2016 =>
            \$v2017\ := \$arr1452_ptr_take\;
            if \$v2017\(0) = '1' then
              \state\ <= q_wait2016;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2014;
            end if;
          when q_wait2022 =>
            \$v2023\ := \$arr1451_ptr_take\;
            if \$v2023\(0) = '1' then
              \state\ <= q_wait2022;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2018\ := "00000000000000000000000000000000";
              \$v2019\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$427_result_after_f\ & "0001" & \$v2018\ & "0001" & \$v2019\;
              \state\ <= pause_setI2020;
            end if;
          when q_wait2028 =>
            \$v2029\ := \$arr1452_ptr_take\;
            if \$v2029\(0) = '1' then
              \state\ <= q_wait2028;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2026;
            end if;
          when q_wait2033 =>
            \$v2034\ := \$arr1451_ptr_take\;
            if \$v2034\(0) = '1' then
              \state\ <= q_wait2033;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2030\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$428_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$427_result_after_f\ & "0010" & \$428_i\ & "0001" & \$v2030\;
              \state\ <= pause_setI2031;
            end if;
          when q_wait2040 =>
            \$v2041\ := \$arr1452_ptr_take\;
            if \$v2041\(0) = '1' then
              \state\ <= q_wait2040;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2038;
            end if;
          when q_wait2056 =>
            \$v2057\ := \$arr1451_ptr_take\;
            if \$v2057\(0) = '1' then
              \state\ <= q_wait2056;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$472\));
              \state\ <= pause_getI2054;
            end if;
          when q_wait2061 =>
            \$v2062\ := \$arr1452_ptr_take\;
            if \$v2062\(0) = '1' then
              \state\ <= q_wait2061;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2059;
            end if;
          when q_wait2065 =>
            \$v2066\ := \$arr1452_ptr_take\;
            if \$v2066\(0) = '1' then
              \state\ <= q_wait2065;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2063;
            end if;
          when q_wait2069 =>
            \$v2070\ := \$arr1451_ptr_take\;
            if \$v2070\(0) = '1' then
              \state\ <= q_wait2069;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$444\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$445\;
              \state\ <= pause_setI2067;
            end if;
          when q_wait2074 =>
            \$v2075\ := \$arr1451_ptr_take\;
            if \$v2075\(0) = '1' then
              \state\ <= q_wait2074;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$452\));
              \state\ <= pause_getI2072;
            end if;
          when q_wait2079 =>
            \$v2080\ := \$arr1452_ptr_take\;
            if \$v2080\(0) = '1' then
              \state\ <= q_wait2079;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2077;
            end if;
          when q_wait2083 =>
            \$v2084\ := \$arr1451_ptr_take\;
            if \$v2084\(0) = '1' then
              \state\ <= q_wait2083;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$458\));
              \state\ <= pause_getI2081;
            end if;
          when q_wait2088 =>
            \$v2089\ := \$arr1452_ptr_take\;
            if \$v2089\(0) = '1' then
              \state\ <= q_wait2088;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2086;
            end if;
          when q_wait2093 =>
            \$v2094\ := \$arr1452_ptr_take\;
            if \$v2094\(0) = '1' then
              \state\ <= q_wait2093;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2091;
            end if;
          when q_wait2101 =>
            \$v2102\ := \$arr1451_ptr_take\;
            if \$v2102\(0) = '1' then
              \state\ <= q_wait2101;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$480\));
              \state\ <= pause_getI2099;
            end if;
          when q_wait2106 =>
            \$v2107\ := \$arr1452_ptr_take\;
            if \$v2107\(0) = '1' then
              \state\ <= q_wait2106;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2104;
            end if;
          when q_wait2110 =>
            \$v2111\ := \$arr1451_ptr_take\;
            if \$v2111\(0) = '1' then
              \state\ <= q_wait2110;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$486\));
              \state\ <= pause_getI2108;
            end if;
          when q_wait2115 =>
            \$v2116\ := \$arr1452_ptr_take\;
            if \$v2116\(0) = '1' then
              \state\ <= q_wait2115;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2113;
            end if;
          when q_wait2124 =>
            \$v2125\ := \$arr1451_ptr_take\;
            if \$v2125\(0) = '1' then
              \state\ <= q_wait2124;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$518\));
              \state\ <= pause_getI2122;
            end if;
          when q_wait2129 =>
            \$v2130\ := \$arr1452_ptr_take\;
            if \$v2130\(0) = '1' then
              \state\ <= q_wait2129;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2127;
            end if;
          when q_wait2133 =>
            \$v2134\ := \$arr1452_ptr_take\;
            if \$v2134\(0) = '1' then
              \state\ <= q_wait2133;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2131;
            end if;
          when q_wait2137 =>
            \$v2138\ := \$arr1451_ptr_take\;
            if \$v2138\(0) = '1' then
              \state\ <= q_wait2137;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$490\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$491\;
              \state\ <= pause_setI2135;
            end if;
          when q_wait2142 =>
            \$v2143\ := \$arr1451_ptr_take\;
            if \$v2143\(0) = '1' then
              \state\ <= q_wait2142;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$498\));
              \state\ <= pause_getI2140;
            end if;
          when q_wait2147 =>
            \$v2148\ := \$arr1452_ptr_take\;
            if \$v2148\(0) = '1' then
              \state\ <= q_wait2147;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2145;
            end if;
          when q_wait2151 =>
            \$v2152\ := \$arr1451_ptr_take\;
            if \$v2152\(0) = '1' then
              \state\ <= q_wait2151;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$504\));
              \state\ <= pause_getI2149;
            end if;
          when q_wait2156 =>
            \$v2157\ := \$arr1452_ptr_take\;
            if \$v2157\(0) = '1' then
              \state\ <= q_wait2156;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2154;
            end if;
          when q_wait2161 =>
            \$v2162\ := \$arr1452_ptr_take\;
            if \$v2162\(0) = '1' then
              \state\ <= q_wait2161;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2159;
            end if;
          when q_wait2169 =>
            \$v2170\ := \$arr1451_ptr_take\;
            if \$v2170\(0) = '1' then
              \state\ <= q_wait2169;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$526\));
              \state\ <= pause_getI2167;
            end if;
          when q_wait2174 =>
            \$v2175\ := \$arr1452_ptr_take\;
            if \$v2175\(0) = '1' then
              \state\ <= q_wait2174;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2172;
            end if;
          when q_wait2178 =>
            \$v2179\ := \$arr1451_ptr_take\;
            if \$v2179\(0) = '1' then
              \state\ <= q_wait2178;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$532\));
              \state\ <= pause_getI2176;
            end if;
          when q_wait2183 =>
            \$v2184\ := \$arr1452_ptr_take\;
            if \$v2184\(0) = '1' then
              \state\ <= q_wait2183;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2181;
            end if;
          when q_wait2187 =>
            \$v2188\ := \$arr1453_ptr_take\;
            if \$v2188\(0) = '1' then
              \state\ <= q_wait2187;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 13;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v108\;
              \state\ <= pause_setI2185;
            end if;
          when q_wait2193 =>
            \$v2194\ := \$arr1452_ptr_take\;
            if \$v2194\(0) = '1' then
              \state\ <= q_wait2193;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2191;
            end if;
          when q_wait2203 =>
            \$v2204\ := \$arr1451_ptr_take\;
            if \$v2204\(0) = '1' then
              \state\ <= q_wait2203;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2198\ := "00000000000000000000000000000000";
              \$v2199\ := "00000000000000000000000000000000";
              \$v2200\ := "00000000000000000000000000000101";
              \$v2195\ := "00000000000000000000000000000000";
              \$v2196\ := "00000000000000000000000000000000";
              \$v2197\ := "00000000000000000000000000000101";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= eclat_if(result & "0001" & \$v2198\ & "0001" & \$v2199\ & "0001" & \$v2200\ & "0001" & \$v2195\ & "0001" & \$v2196\ & "0001" & \$v2197\);
              \state\ <= pause_setI2201;
            end if;
          when q_wait2209 =>
            \$v2210\ := \$arr1452_ptr_take\;
            if \$v2210\(0) = '1' then
              \state\ <= q_wait2209;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2207;
            end if;
          when q_wait2215 =>
            \$v2216\ := \$arr1451_ptr_take\;
            if \$v2216\(0) = '1' then
              \state\ <= q_wait2215;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2211\ := eclat_sub(\$82_i\ & "00000000000000000000000000000001");
              \$v2212\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2211\ & "0010" & \$82_i\ & "0001" & \$v2212\;
              \state\ <= pause_setI2213;
            end if;
          when q_wait2225 =>
            \$v2226\ := \$arr1451_ptr_take\;
            if \$v2226\(0) = '1' then
              \state\ <= q_wait2225;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2220\ := "00000000000000000000000000000000";
              \$v2221\ := "00000000000000000000000000000000";
              \$v2222\ := "00000000000000000000000000000101";
              \$v2217\ := "00000000000000000000000000000000";
              \$v2218\ := "00000000000000000000000000000000";
              \$v2219\ := "00000000000000000000000000000101";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$82_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= eclat_if(result & "0001" & \$v2220\ & "0001" & \$v2221\ & "0001" & \$v2222\ & "0001" & \$v2217\ & "0001" & \$v2218\ & "0001" & \$v2219\);
              \state\ <= pause_setI2223;
            end if;
          when q_wait2232 =>
            \$v2233\ := \$arr1452_ptr_take\;
            if \$v2233\(0) = '1' then
              \state\ <= q_wait2232;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2230;
            end if;
          when q_wait2247 =>
            \$v2248\ := \$arr1451_ptr_take\;
            if \$v2248\(0) = '1' then
              \state\ <= q_wait2247;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$570\));
              \state\ <= pause_getI2245;
            end if;
          when q_wait2252 =>
            \$v2253\ := \$arr1452_ptr_take\;
            if \$v2253\(0) = '1' then
              \state\ <= q_wait2252;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2250;
            end if;
          when q_wait2256 =>
            \$v2257\ := \$arr1452_ptr_take\;
            if \$v2257\(0) = '1' then
              \state\ <= q_wait2256;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2254;
            end if;
          when q_wait2260 =>
            \$v2261\ := \$arr1451_ptr_take\;
            if \$v2261\(0) = '1' then
              \state\ <= q_wait2260;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$542\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$543\;
              \state\ <= pause_setI2258;
            end if;
          when q_wait2265 =>
            \$v2266\ := \$arr1451_ptr_take\;
            if \$v2266\(0) = '1' then
              \state\ <= q_wait2265;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$550\));
              \state\ <= pause_getI2263;
            end if;
          when q_wait2270 =>
            \$v2271\ := \$arr1452_ptr_take\;
            if \$v2271\(0) = '1' then
              \state\ <= q_wait2270;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2268;
            end if;
          when q_wait2274 =>
            \$v2275\ := \$arr1451_ptr_take\;
            if \$v2275\(0) = '1' then
              \state\ <= q_wait2274;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$556\));
              \state\ <= pause_getI2272;
            end if;
          when q_wait2279 =>
            \$v2280\ := \$arr1452_ptr_take\;
            if \$v2280\(0) = '1' then
              \state\ <= q_wait2279;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2277;
            end if;
          when q_wait2284 =>
            \$v2285\ := \$arr1452_ptr_take\;
            if \$v2285\(0) = '1' then
              \state\ <= q_wait2284;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2282;
            end if;
          when q_wait2292 =>
            \$v2293\ := \$arr1451_ptr_take\;
            if \$v2293\(0) = '1' then
              \state\ <= q_wait2292;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$578\));
              \state\ <= pause_getI2290;
            end if;
          when q_wait2297 =>
            \$v2298\ := \$arr1452_ptr_take\;
            if \$v2298\(0) = '1' then
              \state\ <= q_wait2297;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2295;
            end if;
          when q_wait2301 =>
            \$v2302\ := \$arr1451_ptr_take\;
            if \$v2302\(0) = '1' then
              \state\ <= q_wait2301;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$584\));
              \state\ <= pause_getI2299;
            end if;
          when q_wait2306 =>
            \$v2307\ := \$arr1452_ptr_take\;
            if \$v2307\(0) = '1' then
              \state\ <= q_wait2306;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2304;
            end if;
          when q_wait2315 =>
            \$v2316\ := \$arr1451_ptr_take\;
            if \$v2316\(0) = '1' then
              \state\ <= q_wait2315;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$616\));
              \state\ <= pause_getI2313;
            end if;
          when q_wait2320 =>
            \$v2321\ := \$arr1452_ptr_take\;
            if \$v2321\(0) = '1' then
              \state\ <= q_wait2320;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2318;
            end if;
          when q_wait2324 =>
            \$v2325\ := \$arr1452_ptr_take\;
            if \$v2325\(0) = '1' then
              \state\ <= q_wait2324;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2322;
            end if;
          when q_wait2328 =>
            \$v2329\ := \$arr1451_ptr_take\;
            if \$v2329\(0) = '1' then
              \state\ <= q_wait2328;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$588\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$589\;
              \state\ <= pause_setI2326;
            end if;
          when q_wait2333 =>
            \$v2334\ := \$arr1451_ptr_take\;
            if \$v2334\(0) = '1' then
              \state\ <= q_wait2333;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$596\));
              \state\ <= pause_getI2331;
            end if;
          when q_wait2338 =>
            \$v2339\ := \$arr1452_ptr_take\;
            if \$v2339\(0) = '1' then
              \state\ <= q_wait2338;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2336;
            end if;
          when q_wait2342 =>
            \$v2343\ := \$arr1451_ptr_take\;
            if \$v2343\(0) = '1' then
              \state\ <= q_wait2342;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$602\));
              \state\ <= pause_getI2340;
            end if;
          when q_wait2347 =>
            \$v2348\ := \$arr1452_ptr_take\;
            if \$v2348\(0) = '1' then
              \state\ <= q_wait2347;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2345;
            end if;
          when q_wait2352 =>
            \$v2353\ := \$arr1452_ptr_take\;
            if \$v2353\(0) = '1' then
              \state\ <= q_wait2352;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2350;
            end if;
          when q_wait2360 =>
            \$v2361\ := \$arr1451_ptr_take\;
            if \$v2361\(0) = '1' then
              \state\ <= q_wait2360;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$624\));
              \state\ <= pause_getI2358;
            end if;
          when q_wait2365 =>
            \$v2366\ := \$arr1452_ptr_take\;
            if \$v2366\(0) = '1' then
              \state\ <= q_wait2365;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2363;
            end if;
          when q_wait2369 =>
            \$v2370\ := \$arr1451_ptr_take\;
            if \$v2370\(0) = '1' then
              \state\ <= q_wait2369;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$630\));
              \state\ <= pause_getI2367;
            end if;
          when q_wait2374 =>
            \$v2375\ := \$arr1452_ptr_take\;
            if \$v2375\(0) = '1' then
              \state\ <= q_wait2374;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2372;
            end if;
          when q_wait2378 =>
            \$v2379\ := \$arr1453_ptr_take\;
            if \$v2379\(0) = '1' then
              \state\ <= q_wait2378;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 12;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v106\;
              \state\ <= pause_setI2376;
            end if;
          when q_wait2384 =>
            \$v2385\ := \$arr1452_ptr_take\;
            if \$v2385\(0) = '1' then
              \state\ <= q_wait2384;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2382;
            end if;
          when q_wait2394 =>
            \$v2395\ := \$arr1451_ptr_take\;
            if \$v2395\(0) = '1' then
              \state\ <= q_wait2394;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2389\ := "00000000000000000000000000000000";
              \$v2390\ := "00000000000000000000000000000000";
              \$v2391\ := "00000000000000000000000000000101";
              \$v2386\ := "00000000000000000000000000000000";
              \$v2387\ := "00000000000000000000000000000000";
              \$v2388\ := "00000000000000000000000000000101";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2389\ & "0001" & \$v2390\ & "0001" & \$v2391\ & "0001" & \$v2386\ & "0001" & \$v2387\ & "0001" & \$v2388\);
              \state\ <= pause_setI2392;
            end if;
          when q_wait2400 =>
            \$v2401\ := \$arr1452_ptr_take\;
            if \$v2401\(0) = '1' then
              \state\ <= q_wait2400;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2398;
            end if;
          when q_wait2406 =>
            \$v2407\ := \$arr1451_ptr_take\;
            if \$v2407\(0) = '1' then
              \state\ <= q_wait2406;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2402\ := eclat_sub(\$635_i\ & "00000000000000000000000000000001");
              \$v2403\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2402\ & "0010" & \$635_i\ & "0001" & \$v2403\;
              \state\ <= pause_setI2404;
            end if;
          when q_wait2416 =>
            \$v2417\ := \$arr1451_ptr_take\;
            if \$v2417\(0) = '1' then
              \state\ <= q_wait2416;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2411\ := "00000000000000000000000000000000";
              \$v2412\ := "00000000000000000000000000000000";
              \$v2413\ := "00000000000000000000000000000101";
              \$v2408\ := "00000000000000000000000000000000";
              \$v2409\ := "00000000000000000000000000000000";
              \$v2410\ := "00000000000000000000000000000101";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$635_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= eclat_if(\$634_result\ & "0001" & \$v2411\ & "0001" & \$v2412\ & "0001" & \$v2413\ & "0001" & \$v2408\ & "0001" & \$v2409\ & "0001" & \$v2410\);
              \state\ <= pause_setI2414;
            end if;
          when q_wait2423 =>
            \$v2424\ := \$arr1452_ptr_take\;
            if \$v2424\(0) = '1' then
              \state\ <= q_wait2423;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2421;
            end if;
          when q_wait2441 =>
            \$v2442\ := \$arr1451_ptr_take\;
            if \$v2442\(0) = '1' then
              \state\ <= q_wait2441;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$672\));
              \state\ <= pause_getI2439;
            end if;
          when q_wait2446 =>
            \$v2447\ := \$arr1452_ptr_take\;
            if \$v2447\(0) = '1' then
              \state\ <= q_wait2446;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2444;
            end if;
          when q_wait2450 =>
            \$v2451\ := \$arr1452_ptr_take\;
            if \$v2451\(0) = '1' then
              \state\ <= q_wait2450;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2448;
            end if;
          when q_wait2454 =>
            \$v2455\ := \$arr1451_ptr_take\;
            if \$v2455\(0) = '1' then
              \state\ <= q_wait2454;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$644\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$645\;
              \state\ <= pause_setI2452;
            end if;
          when q_wait2459 =>
            \$v2460\ := \$arr1451_ptr_take\;
            if \$v2460\(0) = '1' then
              \state\ <= q_wait2459;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$652\));
              \state\ <= pause_getI2457;
            end if;
          when q_wait2464 =>
            \$v2465\ := \$arr1452_ptr_take\;
            if \$v2465\(0) = '1' then
              \state\ <= q_wait2464;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2462;
            end if;
          when q_wait2468 =>
            \$v2469\ := \$arr1451_ptr_take\;
            if \$v2469\(0) = '1' then
              \state\ <= q_wait2468;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$658\));
              \state\ <= pause_getI2466;
            end if;
          when q_wait2473 =>
            \$v2474\ := \$arr1452_ptr_take\;
            if \$v2474\(0) = '1' then
              \state\ <= q_wait2473;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2471;
            end if;
          when q_wait2478 =>
            \$v2479\ := \$arr1452_ptr_take\;
            if \$v2479\(0) = '1' then
              \state\ <= q_wait2478;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2476;
            end if;
          when q_wait2486 =>
            \$v2487\ := \$arr1451_ptr_take\;
            if \$v2487\(0) = '1' then
              \state\ <= q_wait2486;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$680\));
              \state\ <= pause_getI2484;
            end if;
          when q_wait2491 =>
            \$v2492\ := \$arr1452_ptr_take\;
            if \$v2492\(0) = '1' then
              \state\ <= q_wait2491;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2489;
            end if;
          when q_wait2495 =>
            \$v2496\ := \$arr1451_ptr_take\;
            if \$v2496\(0) = '1' then
              \state\ <= q_wait2495;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$686\));
              \state\ <= pause_getI2493;
            end if;
          when q_wait2500 =>
            \$v2501\ := \$arr1452_ptr_take\;
            if \$v2501\(0) = '1' then
              \state\ <= q_wait2500;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2498;
            end if;
          when q_wait2509 =>
            \$v2510\ := \$arr1451_ptr_take\;
            if \$v2510\(0) = '1' then
              \state\ <= q_wait2509;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$718\));
              \state\ <= pause_getI2507;
            end if;
          when q_wait2514 =>
            \$v2515\ := \$arr1452_ptr_take\;
            if \$v2515\(0) = '1' then
              \state\ <= q_wait2514;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2512;
            end if;
          when q_wait2518 =>
            \$v2519\ := \$arr1452_ptr_take\;
            if \$v2519\(0) = '1' then
              \state\ <= q_wait2518;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2516;
            end if;
          when q_wait2522 =>
            \$v2523\ := \$arr1451_ptr_take\;
            if \$v2523\(0) = '1' then
              \state\ <= q_wait2522;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$690\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$691\;
              \state\ <= pause_setI2520;
            end if;
          when q_wait2527 =>
            \$v2528\ := \$arr1451_ptr_take\;
            if \$v2528\(0) = '1' then
              \state\ <= q_wait2527;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$698\));
              \state\ <= pause_getI2525;
            end if;
          when q_wait2532 =>
            \$v2533\ := \$arr1452_ptr_take\;
            if \$v2533\(0) = '1' then
              \state\ <= q_wait2532;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2530;
            end if;
          when q_wait2536 =>
            \$v2537\ := \$arr1451_ptr_take\;
            if \$v2537\(0) = '1' then
              \state\ <= q_wait2536;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$704\));
              \state\ <= pause_getI2534;
            end if;
          when q_wait2541 =>
            \$v2542\ := \$arr1452_ptr_take\;
            if \$v2542\(0) = '1' then
              \state\ <= q_wait2541;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2539;
            end if;
          when q_wait2546 =>
            \$v2547\ := \$arr1452_ptr_take\;
            if \$v2547\(0) = '1' then
              \state\ <= q_wait2546;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2544;
            end if;
          when q_wait2554 =>
            \$v2555\ := \$arr1451_ptr_take\;
            if \$v2555\(0) = '1' then
              \state\ <= q_wait2554;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$726\));
              \state\ <= pause_getI2552;
            end if;
          when q_wait2559 =>
            \$v2560\ := \$arr1452_ptr_take\;
            if \$v2560\(0) = '1' then
              \state\ <= q_wait2559;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2557;
            end if;
          when q_wait2563 =>
            \$v2564\ := \$arr1451_ptr_take\;
            if \$v2564\(0) = '1' then
              \state\ <= q_wait2563;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$732\));
              \state\ <= pause_getI2561;
            end if;
          when q_wait2568 =>
            \$v2569\ := \$arr1452_ptr_take\;
            if \$v2569\(0) = '1' then
              \state\ <= q_wait2568;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2566;
            end if;
          when q_wait2572 =>
            \$v2573\ := \$arr1453_ptr_take\;
            if \$v2573\(0) = '1' then
              \state\ <= q_wait2572;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 11;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v104\;
              \state\ <= pause_setI2570;
            end if;
          when q_wait2578 =>
            \$v2579\ := \$arr1452_ptr_take\;
            if \$v2579\(0) = '1' then
              \state\ <= q_wait2578;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2576;
            end if;
          when q_wait2582 =>
            \$v2583\ := \$arr1451_ptr_take\;
            if \$v2583\(0) = '1' then
              \state\ <= q_wait2582;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
              \state\ <= pause_setI2580;
            end if;
          when q_wait2588 =>
            \$v2589\ := \$arr1452_ptr_take\;
            if \$v2589\(0) = '1' then
              \state\ <= q_wait2588;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2586;
            end if;
          when q_wait2594 =>
            \$v2595\ := \$arr1451_ptr_take\;
            if \$v2595\(0) = '1' then
              \state\ <= q_wait2594;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2590\ := eclat_sub(\$734_i\ & "00000000000000000000000000000001");
              \$v2591\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2590\ & "0010" & \$734_i\ & "0001" & \$v2591\;
              \state\ <= pause_setI2592;
            end if;
          when q_wait2598 =>
            \$v2599\ := \$arr1451_ptr_take\;
            if \$v2599\(0) = '1' then
              \state\ <= q_wait2598;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$734_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$56_y\(0 to 35) & \$56_y\(36 to 71) & \$55_x\;
              \state\ <= pause_setI2596;
            end if;
          when q_wait2605 =>
            \$v2606\ := \$arr1452_ptr_take\;
            if \$v2606\(0) = '1' then
              \state\ <= q_wait2605;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2603;
            end if;
          when q_wait2610 =>
            \$v2611\ := \$arr1451_ptr_take\;
            if \$v2611\(0) = '1' then
              \state\ <= q_wait2610;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$135_i\));
              \state\ <= pause_getI2608;
            end if;
          when q_wait2621 =>
            \$v2622\ := \$arr1451_ptr_take\;
            if \$v2622\(0) = '1' then
              \state\ <= q_wait2621;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$777\));
              \state\ <= pause_getI2619;
            end if;
          when q_wait2626 =>
            \$v2627\ := \$arr1452_ptr_take\;
            if \$v2627\(0) = '1' then
              \state\ <= q_wait2626;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2624;
            end if;
          when q_wait2630 =>
            \$v2631\ := \$arr1452_ptr_take\;
            if \$v2631\(0) = '1' then
              \state\ <= q_wait2630;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2628;
            end if;
          when q_wait2634 =>
            \$v2635\ := \$arr1451_ptr_take\;
            if \$v2635\(0) = '1' then
              \state\ <= q_wait2634;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$749\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$750\;
              \state\ <= pause_setI2632;
            end if;
          when q_wait2639 =>
            \$v2640\ := \$arr1451_ptr_take\;
            if \$v2640\(0) = '1' then
              \state\ <= q_wait2639;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$757\));
              \state\ <= pause_getI2637;
            end if;
          when q_wait2644 =>
            \$v2645\ := \$arr1452_ptr_take\;
            if \$v2645\(0) = '1' then
              \state\ <= q_wait2644;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2642;
            end if;
          when q_wait2648 =>
            \$v2649\ := \$arr1451_ptr_take\;
            if \$v2649\(0) = '1' then
              \state\ <= q_wait2648;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$763\));
              \state\ <= pause_getI2646;
            end if;
          when q_wait2653 =>
            \$v2654\ := \$arr1452_ptr_take\;
            if \$v2654\(0) = '1' then
              \state\ <= q_wait2653;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2651;
            end if;
          when q_wait2658 =>
            \$v2659\ := \$arr1452_ptr_take\;
            if \$v2659\(0) = '1' then
              \state\ <= q_wait2658;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2656;
            end if;
          when q_wait2666 =>
            \$v2667\ := \$arr1451_ptr_take\;
            if \$v2667\(0) = '1' then
              \state\ <= q_wait2666;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$785\));
              \state\ <= pause_getI2664;
            end if;
          when q_wait2671 =>
            \$v2672\ := \$arr1452_ptr_take\;
            if \$v2672\(0) = '1' then
              \state\ <= q_wait2671;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2669;
            end if;
          when q_wait2675 =>
            \$v2676\ := \$arr1451_ptr_take\;
            if \$v2676\(0) = '1' then
              \state\ <= q_wait2675;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$791\));
              \state\ <= pause_getI2673;
            end if;
          when q_wait2680 =>
            \$v2681\ := \$arr1452_ptr_take\;
            if \$v2681\(0) = '1' then
              \state\ <= q_wait2680;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2678;
            end if;
          when q_wait2689 =>
            \$v2690\ := \$arr1451_ptr_take\;
            if \$v2690\(0) = '1' then
              \state\ <= q_wait2689;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$823\));
              \state\ <= pause_getI2687;
            end if;
          when q_wait2694 =>
            \$v2695\ := \$arr1452_ptr_take\;
            if \$v2695\(0) = '1' then
              \state\ <= q_wait2694;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2692;
            end if;
          when q_wait2698 =>
            \$v2699\ := \$arr1452_ptr_take\;
            if \$v2699\(0) = '1' then
              \state\ <= q_wait2698;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2696;
            end if;
          when q_wait2702 =>
            \$v2703\ := \$arr1451_ptr_take\;
            if \$v2703\(0) = '1' then
              \state\ <= q_wait2702;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$795\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$796\;
              \state\ <= pause_setI2700;
            end if;
          when q_wait2707 =>
            \$v2708\ := \$arr1451_ptr_take\;
            if \$v2708\(0) = '1' then
              \state\ <= q_wait2707;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$803\));
              \state\ <= pause_getI2705;
            end if;
          when q_wait2712 =>
            \$v2713\ := \$arr1452_ptr_take\;
            if \$v2713\(0) = '1' then
              \state\ <= q_wait2712;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2710;
            end if;
          when q_wait2716 =>
            \$v2717\ := \$arr1451_ptr_take\;
            if \$v2717\(0) = '1' then
              \state\ <= q_wait2716;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$809\));
              \state\ <= pause_getI2714;
            end if;
          when q_wait2721 =>
            \$v2722\ := \$arr1452_ptr_take\;
            if \$v2722\(0) = '1' then
              \state\ <= q_wait2721;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2719;
            end if;
          when q_wait2726 =>
            \$v2727\ := \$arr1452_ptr_take\;
            if \$v2727\(0) = '1' then
              \state\ <= q_wait2726;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2724;
            end if;
          when q_wait2734 =>
            \$v2735\ := \$arr1451_ptr_take\;
            if \$v2735\(0) = '1' then
              \state\ <= q_wait2734;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$831\));
              \state\ <= pause_getI2732;
            end if;
          when q_wait2739 =>
            \$v2740\ := \$arr1452_ptr_take\;
            if \$v2740\(0) = '1' then
              \state\ <= q_wait2739;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2737;
            end if;
          when q_wait2743 =>
            \$v2744\ := \$arr1451_ptr_take\;
            if \$v2744\(0) = '1' then
              \state\ <= q_wait2743;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$837\));
              \state\ <= pause_getI2741;
            end if;
          when q_wait2748 =>
            \$v2749\ := \$arr1452_ptr_take\;
            if \$v2749\(0) = '1' then
              \state\ <= q_wait2748;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2746;
            end if;
          when q_wait2752 =>
            \$v2753\ := \$arr1453_ptr_take\;
            if \$v2753\(0) = '1' then
              \state\ <= q_wait2752;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 10;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v102\;
              \state\ <= pause_setI2750;
            end if;
          when q_wait2758 =>
            \$v2759\ := \$arr1452_ptr_take\;
            if \$v2759\(0) = '1' then
              \state\ <= q_wait2758;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2756;
            end if;
          when q_wait2762 =>
            \$v2763\ := \$arr1451_ptr_take\;
            if \$v2763\(0) = '1' then
              \state\ <= q_wait2762;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
              \state\ <= pause_setI2760;
            end if;
          when q_wait2768 =>
            \$v2769\ := \$arr1452_ptr_take\;
            if \$v2769\(0) = '1' then
              \state\ <= q_wait2768;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2766;
            end if;
          when q_wait2774 =>
            \$v2775\ := \$arr1451_ptr_take\;
            if \$v2775\(0) = '1' then
              \state\ <= q_wait2774;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2770\ := eclat_sub(\$841_i\ & "00000000000000000000000000000001");
              \$v2771\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2770\ & "0010" & \$841_i\ & "0001" & \$v2771\;
              \state\ <= pause_setI2772;
            end if;
          when q_wait2778 =>
            \$v2779\ := \$arr1451_ptr_take\;
            if \$v2779\(0) = '1' then
              \state\ <= q_wait2778;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$841_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$840_y\(0 to 35) & \$839_x\ & \$840_y\(72 to 107);
              \state\ <= pause_setI2776;
            end if;
          when q_wait2785 =>
            \$v2786\ := \$arr1452_ptr_take\;
            if \$v2786\(0) = '1' then
              \state\ <= q_wait2785;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2783;
            end if;
          when q_wait2790 =>
            \$v2791\ := \$arr1451_ptr_take\;
            if \$v2791\(0) = '1' then
              \state\ <= q_wait2790;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$852_i\));
              \state\ <= pause_getI2788;
            end if;
          when q_wait2801 =>
            \$v2802\ := \$arr1451_ptr_take\;
            if \$v2802\(0) = '1' then
              \state\ <= q_wait2801;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$886\));
              \state\ <= pause_getI2799;
            end if;
          when q_wait2806 =>
            \$v2807\ := \$arr1452_ptr_take\;
            if \$v2807\(0) = '1' then
              \state\ <= q_wait2806;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2804;
            end if;
          when q_wait2810 =>
            \$v2811\ := \$arr1452_ptr_take\;
            if \$v2811\(0) = '1' then
              \state\ <= q_wait2810;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2808;
            end if;
          when q_wait2814 =>
            \$v2815\ := \$arr1451_ptr_take\;
            if \$v2815\(0) = '1' then
              \state\ <= q_wait2814;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$858\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$859\;
              \state\ <= pause_setI2812;
            end if;
          when q_wait2819 =>
            \$v2820\ := \$arr1451_ptr_take\;
            if \$v2820\(0) = '1' then
              \state\ <= q_wait2819;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$866\));
              \state\ <= pause_getI2817;
            end if;
          when q_wait2824 =>
            \$v2825\ := \$arr1452_ptr_take\;
            if \$v2825\(0) = '1' then
              \state\ <= q_wait2824;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2822;
            end if;
          when q_wait2828 =>
            \$v2829\ := \$arr1451_ptr_take\;
            if \$v2829\(0) = '1' then
              \state\ <= q_wait2828;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$872\));
              \state\ <= pause_getI2826;
            end if;
          when q_wait2833 =>
            \$v2834\ := \$arr1452_ptr_take\;
            if \$v2834\(0) = '1' then
              \state\ <= q_wait2833;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2831;
            end if;
          when q_wait2838 =>
            \$v2839\ := \$arr1452_ptr_take\;
            if \$v2839\(0) = '1' then
              \state\ <= q_wait2838;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2836;
            end if;
          when q_wait2846 =>
            \$v2847\ := \$arr1451_ptr_take\;
            if \$v2847\(0) = '1' then
              \state\ <= q_wait2846;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$894\));
              \state\ <= pause_getI2844;
            end if;
          when q_wait2851 =>
            \$v2852\ := \$arr1452_ptr_take\;
            if \$v2852\(0) = '1' then
              \state\ <= q_wait2851;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2849;
            end if;
          when q_wait2855 =>
            \$v2856\ := \$arr1451_ptr_take\;
            if \$v2856\(0) = '1' then
              \state\ <= q_wait2855;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$900\));
              \state\ <= pause_getI2853;
            end if;
          when q_wait2860 =>
            \$v2861\ := \$arr1452_ptr_take\;
            if \$v2861\(0) = '1' then
              \state\ <= q_wait2860;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2858;
            end if;
          when q_wait2869 =>
            \$v2870\ := \$arr1451_ptr_take\;
            if \$v2870\(0) = '1' then
              \state\ <= q_wait2869;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$932\));
              \state\ <= pause_getI2867;
            end if;
          when q_wait2874 =>
            \$v2875\ := \$arr1452_ptr_take\;
            if \$v2875\(0) = '1' then
              \state\ <= q_wait2874;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2872;
            end if;
          when q_wait2878 =>
            \$v2879\ := \$arr1452_ptr_take\;
            if \$v2879\(0) = '1' then
              \state\ <= q_wait2878;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2876;
            end if;
          when q_wait2882 =>
            \$v2883\ := \$arr1451_ptr_take\;
            if \$v2883\(0) = '1' then
              \state\ <= q_wait2882;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$904\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$905\;
              \state\ <= pause_setI2880;
            end if;
          when q_wait2887 =>
            \$v2888\ := \$arr1451_ptr_take\;
            if \$v2888\(0) = '1' then
              \state\ <= q_wait2887;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$912\));
              \state\ <= pause_getI2885;
            end if;
          when q_wait2892 =>
            \$v2893\ := \$arr1452_ptr_take\;
            if \$v2893\(0) = '1' then
              \state\ <= q_wait2892;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2890;
            end if;
          when q_wait2896 =>
            \$v2897\ := \$arr1451_ptr_take\;
            if \$v2897\(0) = '1' then
              \state\ <= q_wait2896;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$918\));
              \state\ <= pause_getI2894;
            end if;
          when q_wait2901 =>
            \$v2902\ := \$arr1452_ptr_take\;
            if \$v2902\(0) = '1' then
              \state\ <= q_wait2901;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2899;
            end if;
          when q_wait2906 =>
            \$v2907\ := \$arr1452_ptr_take\;
            if \$v2907\(0) = '1' then
              \state\ <= q_wait2906;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2904;
            end if;
          when q_wait2914 =>
            \$v2915\ := \$arr1451_ptr_take\;
            if \$v2915\(0) = '1' then
              \state\ <= q_wait2914;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$940\));
              \state\ <= pause_getI2912;
            end if;
          when q_wait2919 =>
            \$v2920\ := \$arr1452_ptr_take\;
            if \$v2920\(0) = '1' then
              \state\ <= q_wait2919;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2917;
            end if;
          when q_wait2923 =>
            \$v2924\ := \$arr1451_ptr_take\;
            if \$v2924\(0) = '1' then
              \state\ <= q_wait2923;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$946\));
              \state\ <= pause_getI2921;
            end if;
          when q_wait2928 =>
            \$v2929\ := \$arr1452_ptr_take\;
            if \$v2929\(0) = '1' then
              \state\ <= q_wait2928;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2926;
            end if;
          when q_wait2932 =>
            \$v2933\ := \$arr1453_ptr_take\;
            if \$v2933\(0) = '1' then
              \state\ <= q_wait2932;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 9;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v100\;
              \state\ <= pause_setI2930;
            end if;
          when q_wait2938 =>
            \$v2939\ := \$arr1452_ptr_take\;
            if \$v2939\(0) = '1' then
              \state\ <= q_wait2938;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2936;
            end if;
          when q_wait2942 =>
            \$v2943\ := \$arr1451_ptr_take\;
            if \$v2943\(0) = '1' then
              \state\ <= q_wait2942;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
              \state\ <= pause_setI2940;
            end if;
          when q_wait2948 =>
            \$v2949\ := \$arr1452_ptr_take\;
            if \$v2949\(0) = '1' then
              \state\ <= q_wait2948;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2946;
            end if;
          when q_wait2954 =>
            \$v2955\ := \$arr1451_ptr_take\;
            if \$v2955\(0) = '1' then
              \state\ <= q_wait2954;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v2950\ := eclat_sub(\$950_i\ & "00000000000000000000000000000001");
              \$v2951\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v2950\ & "0010" & \$950_i\ & "0001" & \$v2951\;
              \state\ <= pause_setI2952;
            end if;
          when q_wait2958 =>
            \$v2959\ := \$arr1451_ptr_take\;
            if \$v2959\(0) = '1' then
              \state\ <= q_wait2958;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$950_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$948_x\ & \$949_y\(36 to 71) & \$949_y\(72 to 107);
              \state\ <= pause_setI2956;
            end if;
          when q_wait2965 =>
            \$v2966\ := \$arr1452_ptr_take\;
            if \$v2966\(0) = '1' then
              \state\ <= q_wait2965;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2963;
            end if;
          when q_wait2970 =>
            \$v2971\ := \$arr1451_ptr_take\;
            if \$v2971\(0) = '1' then
              \state\ <= q_wait2970;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$961_i\));
              \state\ <= pause_getI2968;
            end if;
          when q_wait2981 =>
            \$v2982\ := \$arr1451_ptr_take\;
            if \$v2982\(0) = '1' then
              \state\ <= q_wait2981;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$995\));
              \state\ <= pause_getI2979;
            end if;
          when q_wait2986 =>
            \$v2987\ := \$arr1452_ptr_take\;
            if \$v2987\(0) = '1' then
              \state\ <= q_wait2986;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2984;
            end if;
          when q_wait2990 =>
            \$v2991\ := \$arr1452_ptr_take\;
            if \$v2991\(0) = '1' then
              \state\ <= q_wait2990;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI2988;
            end if;
          when q_wait2994 =>
            \$v2995\ := \$arr1451_ptr_take\;
            if \$v2995\(0) = '1' then
              \state\ <= q_wait2994;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$967\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$968\;
              \state\ <= pause_setI2992;
            end if;
          when q_wait2999 =>
            \$v3000\ := \$arr1451_ptr_take\;
            if \$v3000\(0) = '1' then
              \state\ <= q_wait2999;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$975\));
              \state\ <= pause_getI2997;
            end if;
          when q_wait3004 =>
            \$v3005\ := \$arr1452_ptr_take\;
            if \$v3005\(0) = '1' then
              \state\ <= q_wait3004;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3002;
            end if;
          when q_wait3008 =>
            \$v3009\ := \$arr1451_ptr_take\;
            if \$v3009\(0) = '1' then
              \state\ <= q_wait3008;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$981\));
              \state\ <= pause_getI3006;
            end if;
          when q_wait3013 =>
            \$v3014\ := \$arr1452_ptr_take\;
            if \$v3014\(0) = '1' then
              \state\ <= q_wait3013;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3011;
            end if;
          when q_wait3018 =>
            \$v3019\ := \$arr1452_ptr_take\;
            if \$v3019\(0) = '1' then
              \state\ <= q_wait3018;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3016;
            end if;
          when q_wait3026 =>
            \$v3027\ := \$arr1451_ptr_take\;
            if \$v3027\(0) = '1' then
              \state\ <= q_wait3026;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1003\));
              \state\ <= pause_getI3024;
            end if;
          when q_wait3031 =>
            \$v3032\ := \$arr1452_ptr_take\;
            if \$v3032\(0) = '1' then
              \state\ <= q_wait3031;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3029;
            end if;
          when q_wait3035 =>
            \$v3036\ := \$arr1451_ptr_take\;
            if \$v3036\(0) = '1' then
              \state\ <= q_wait3035;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1009\));
              \state\ <= pause_getI3033;
            end if;
          when q_wait3040 =>
            \$v3041\ := \$arr1452_ptr_take\;
            if \$v3041\(0) = '1' then
              \state\ <= q_wait3040;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3038;
            end if;
          when q_wait3049 =>
            \$v3050\ := \$arr1451_ptr_take\;
            if \$v3050\(0) = '1' then
              \state\ <= q_wait3049;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1041\));
              \state\ <= pause_getI3047;
            end if;
          when q_wait3054 =>
            \$v3055\ := \$arr1452_ptr_take\;
            if \$v3055\(0) = '1' then
              \state\ <= q_wait3054;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3052;
            end if;
          when q_wait3058 =>
            \$v3059\ := \$arr1452_ptr_take\;
            if \$v3059\(0) = '1' then
              \state\ <= q_wait3058;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3056;
            end if;
          when q_wait3062 =>
            \$v3063\ := \$arr1451_ptr_take\;
            if \$v3063\(0) = '1' then
              \state\ <= q_wait3062;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1013\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1014\;
              \state\ <= pause_setI3060;
            end if;
          when q_wait3067 =>
            \$v3068\ := \$arr1451_ptr_take\;
            if \$v3068\(0) = '1' then
              \state\ <= q_wait3067;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1021\));
              \state\ <= pause_getI3065;
            end if;
          when q_wait3072 =>
            \$v3073\ := \$arr1452_ptr_take\;
            if \$v3073\(0) = '1' then
              \state\ <= q_wait3072;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3070;
            end if;
          when q_wait3076 =>
            \$v3077\ := \$arr1451_ptr_take\;
            if \$v3077\(0) = '1' then
              \state\ <= q_wait3076;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1027\));
              \state\ <= pause_getI3074;
            end if;
          when q_wait3081 =>
            \$v3082\ := \$arr1452_ptr_take\;
            if \$v3082\(0) = '1' then
              \state\ <= q_wait3081;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3079;
            end if;
          when q_wait3086 =>
            \$v3087\ := \$arr1452_ptr_take\;
            if \$v3087\(0) = '1' then
              \state\ <= q_wait3086;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3084;
            end if;
          when q_wait3094 =>
            \$v3095\ := \$arr1451_ptr_take\;
            if \$v3095\(0) = '1' then
              \state\ <= q_wait3094;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1049\));
              \state\ <= pause_getI3092;
            end if;
          when q_wait3099 =>
            \$v3100\ := \$arr1452_ptr_take\;
            if \$v3100\(0) = '1' then
              \state\ <= q_wait3099;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3097;
            end if;
          when q_wait3103 =>
            \$v3104\ := \$arr1451_ptr_take\;
            if \$v3104\(0) = '1' then
              \state\ <= q_wait3103;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1055\));
              \state\ <= pause_getI3101;
            end if;
          when q_wait3108 =>
            \$v3109\ := \$arr1452_ptr_take\;
            if \$v3109\(0) = '1' then
              \state\ <= q_wait3108;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3106;
            end if;
          when q_wait3112 =>
            \$v3113\ := \$arr1453_ptr_take\;
            if \$v3113\(0) = '1' then
              \state\ <= q_wait3112;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 8;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v98\;
              \state\ <= pause_setI3110;
            end if;
          when q_wait3119 =>
            \$v3120\ := \$arr1452_ptr_take\;
            if \$v3120\(0) = '1' then
              \state\ <= q_wait3119;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3117;
            end if;
          when q_wait3123 =>
            \$v3124\ := \$arr1452_ptr_take\;
            if \$v3124\(0) = '1' then
              \state\ <= q_wait3123;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3121;
            end if;
          when q_wait3129 =>
            \$v3130\ := \$arr1451_ptr_take\;
            if \$v3130\(0) = '1' then
              \state\ <= q_wait3129;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3125\ := "00000000000000000000000000000000";
              \$v3126\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$58_result\(72 to 107) & "0001" & \$v3125\ & "0001" & \$v3126\;
              \state\ <= pause_setI3127;
            end if;
          when q_wait3135 =>
            \$v3136\ := \$arr1452_ptr_take\;
            if \$v3136\(0) = '1' then
              \state\ <= q_wait3135;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3133;
            end if;
          when q_wait3140 =>
            \$v3141\ := \$arr1451_ptr_take\;
            if \$v3141\(0) = '1' then
              \state\ <= q_wait3140;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3137\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1057_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$58_result\(72 to 107) & "0010" & \$1057_i\ & "0001" & \$v3137\;
              \state\ <= pause_setI3138;
            end if;
          when q_wait3147 =>
            \$v3148\ := \$arr1452_ptr_take\;
            if \$v3148\(0) = '1' then
              \state\ <= q_wait3147;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3145;
            end if;
          when q_wait3152 =>
            \$v3153\ := \$arr1451_ptr_take\;
            if \$v3153\(0) = '1' then
              \state\ <= q_wait3152;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1075_i\));
              \state\ <= pause_getI3150;
            end if;
          when q_wait3163 =>
            \$v3164\ := \$arr1451_ptr_take\;
            if \$v3164\(0) = '1' then
              \state\ <= q_wait3163;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1109\));
              \state\ <= pause_getI3161;
            end if;
          when q_wait3168 =>
            \$v3169\ := \$arr1452_ptr_take\;
            if \$v3169\(0) = '1' then
              \state\ <= q_wait3168;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3166;
            end if;
          when q_wait3172 =>
            \$v3173\ := \$arr1452_ptr_take\;
            if \$v3173\(0) = '1' then
              \state\ <= q_wait3172;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3170;
            end if;
          when q_wait3176 =>
            \$v3177\ := \$arr1451_ptr_take\;
            if \$v3177\(0) = '1' then
              \state\ <= q_wait3176;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1081\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1082\;
              \state\ <= pause_setI3174;
            end if;
          when q_wait3181 =>
            \$v3182\ := \$arr1451_ptr_take\;
            if \$v3182\(0) = '1' then
              \state\ <= q_wait3181;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1089\));
              \state\ <= pause_getI3179;
            end if;
          when q_wait3186 =>
            \$v3187\ := \$arr1452_ptr_take\;
            if \$v3187\(0) = '1' then
              \state\ <= q_wait3186;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3184;
            end if;
          when q_wait3190 =>
            \$v3191\ := \$arr1451_ptr_take\;
            if \$v3191\(0) = '1' then
              \state\ <= q_wait3190;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1095\));
              \state\ <= pause_getI3188;
            end if;
          when q_wait3195 =>
            \$v3196\ := \$arr1452_ptr_take\;
            if \$v3196\(0) = '1' then
              \state\ <= q_wait3195;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3193;
            end if;
          when q_wait3200 =>
            \$v3201\ := \$arr1452_ptr_take\;
            if \$v3201\(0) = '1' then
              \state\ <= q_wait3200;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3198;
            end if;
          when q_wait3208 =>
            \$v3209\ := \$arr1451_ptr_take\;
            if \$v3209\(0) = '1' then
              \state\ <= q_wait3208;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1117\));
              \state\ <= pause_getI3206;
            end if;
          when q_wait3213 =>
            \$v3214\ := \$arr1452_ptr_take\;
            if \$v3214\(0) = '1' then
              \state\ <= q_wait3213;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3211;
            end if;
          when q_wait3217 =>
            \$v3218\ := \$arr1451_ptr_take\;
            if \$v3218\(0) = '1' then
              \state\ <= q_wait3217;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1123\));
              \state\ <= pause_getI3215;
            end if;
          when q_wait3222 =>
            \$v3223\ := \$arr1452_ptr_take\;
            if \$v3223\(0) = '1' then
              \state\ <= q_wait3222;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3220;
            end if;
          when q_wait3226 =>
            \$v3227\ := \$arr1453_ptr_take\;
            if \$v3227\(0) = '1' then
              \state\ <= q_wait3226;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 7;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v97\;
              \state\ <= pause_setI3224;
            end if;
          when q_wait3233 =>
            \$v3234\ := \$arr1452_ptr_take\;
            if \$v3234\(0) = '1' then
              \state\ <= q_wait3233;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3231;
            end if;
          when q_wait3237 =>
            \$v3238\ := \$arr1452_ptr_take\;
            if \$v3238\(0) = '1' then
              \state\ <= q_wait3237;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3235;
            end if;
          when q_wait3243 =>
            \$v3244\ := \$arr1451_ptr_take\;
            if \$v3244\(0) = '1' then
              \state\ <= q_wait3243;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3239\ := "00000000000000000000000000000000";
              \$v3240\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1125_result\(36 to 71) & "0001" & \$v3239\ & "0001" & \$v3240\;
              \state\ <= pause_setI3241;
            end if;
          when q_wait3249 =>
            \$v3250\ := \$arr1452_ptr_take\;
            if \$v3250\(0) = '1' then
              \state\ <= q_wait3249;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3247;
            end if;
          when q_wait3254 =>
            \$v3255\ := \$arr1451_ptr_take\;
            if \$v3255\(0) = '1' then
              \state\ <= q_wait3254;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3251\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1126_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1125_result\(36 to 71) & "0010" & \$1126_i\ & "0001" & \$v3251\;
              \state\ <= pause_setI3252;
            end if;
          when q_wait3261 =>
            \$v3262\ := \$arr1452_ptr_take\;
            if \$v3262\(0) = '1' then
              \state\ <= q_wait3261;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3259;
            end if;
          when q_wait3266 =>
            \$v3267\ := \$arr1451_ptr_take\;
            if \$v3267\(0) = '1' then
              \state\ <= q_wait3266;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1144_i\));
              \state\ <= pause_getI3264;
            end if;
          when q_wait3277 =>
            \$v3278\ := \$arr1451_ptr_take\;
            if \$v3278\(0) = '1' then
              \state\ <= q_wait3277;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1178\));
              \state\ <= pause_getI3275;
            end if;
          when q_wait3282 =>
            \$v3283\ := \$arr1452_ptr_take\;
            if \$v3283\(0) = '1' then
              \state\ <= q_wait3282;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3280;
            end if;
          when q_wait3286 =>
            \$v3287\ := \$arr1452_ptr_take\;
            if \$v3287\(0) = '1' then
              \state\ <= q_wait3286;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3284;
            end if;
          when q_wait3290 =>
            \$v3291\ := \$arr1451_ptr_take\;
            if \$v3291\(0) = '1' then
              \state\ <= q_wait3290;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1150\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1151\;
              \state\ <= pause_setI3288;
            end if;
          when q_wait3295 =>
            \$v3296\ := \$arr1451_ptr_take\;
            if \$v3296\(0) = '1' then
              \state\ <= q_wait3295;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1158\));
              \state\ <= pause_getI3293;
            end if;
          when q_wait3300 =>
            \$v3301\ := \$arr1452_ptr_take\;
            if \$v3301\(0) = '1' then
              \state\ <= q_wait3300;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3298;
            end if;
          when q_wait3304 =>
            \$v3305\ := \$arr1451_ptr_take\;
            if \$v3305\(0) = '1' then
              \state\ <= q_wait3304;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1164\));
              \state\ <= pause_getI3302;
            end if;
          when q_wait3309 =>
            \$v3310\ := \$arr1452_ptr_take\;
            if \$v3310\(0) = '1' then
              \state\ <= q_wait3309;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3307;
            end if;
          when q_wait3314 =>
            \$v3315\ := \$arr1452_ptr_take\;
            if \$v3315\(0) = '1' then
              \state\ <= q_wait3314;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3312;
            end if;
          when q_wait3322 =>
            \$v3323\ := \$arr1451_ptr_take\;
            if \$v3323\(0) = '1' then
              \state\ <= q_wait3322;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1186\));
              \state\ <= pause_getI3320;
            end if;
          when q_wait3327 =>
            \$v3328\ := \$arr1452_ptr_take\;
            if \$v3328\(0) = '1' then
              \state\ <= q_wait3327;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3325;
            end if;
          when q_wait3331 =>
            \$v3332\ := \$arr1451_ptr_take\;
            if \$v3332\(0) = '1' then
              \state\ <= q_wait3331;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1192\));
              \state\ <= pause_getI3329;
            end if;
          when q_wait3336 =>
            \$v3337\ := \$arr1452_ptr_take\;
            if \$v3337\(0) = '1' then
              \state\ <= q_wait3336;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3334;
            end if;
          when q_wait3340 =>
            \$v3341\ := \$arr1453_ptr_take\;
            if \$v3341\(0) = '1' then
              \state\ <= q_wait3340;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 6;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v96\;
              \state\ <= pause_setI3338;
            end if;
          when q_wait3347 =>
            \$v3348\ := \$arr1452_ptr_take\;
            if \$v3348\(0) = '1' then
              \state\ <= q_wait3347;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3345;
            end if;
          when q_wait3351 =>
            \$v3352\ := \$arr1452_ptr_take\;
            if \$v3352\(0) = '1' then
              \state\ <= q_wait3351;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3349;
            end if;
          when q_wait3357 =>
            \$v3358\ := \$arr1451_ptr_take\;
            if \$v3358\(0) = '1' then
              \state\ <= q_wait3357;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3353\ := "00000000000000000000000000000000";
              \$v3354\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1194_result\(0 to 35) & "0001" & \$v3353\ & "0001" & \$v3354\;
              \state\ <= pause_setI3355;
            end if;
          when q_wait3363 =>
            \$v3364\ := \$arr1452_ptr_take\;
            if \$v3364\(0) = '1' then
              \state\ <= q_wait3363;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3361;
            end if;
          when q_wait3368 =>
            \$v3369\ := \$arr1451_ptr_take\;
            if \$v3369\(0) = '1' then
              \state\ <= q_wait3368;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3365\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1195_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1194_result\(0 to 35) & "0010" & \$1195_i\ & "0001" & \$v3365\;
              \state\ <= pause_setI3366;
            end if;
          when q_wait3375 =>
            \$v3376\ := \$arr1452_ptr_take\;
            if \$v3376\(0) = '1' then
              \state\ <= q_wait3375;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3373;
            end if;
          when q_wait3380 =>
            \$v3381\ := \$arr1451_ptr_take\;
            if \$v3381\(0) = '1' then
              \state\ <= q_wait3380;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1213_i\));
              \state\ <= pause_getI3378;
            end if;
          when q_wait3391 =>
            \$v3392\ := \$arr1451_ptr_take\;
            if \$v3392\(0) = '1' then
              \state\ <= q_wait3391;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1247\));
              \state\ <= pause_getI3389;
            end if;
          when q_wait3396 =>
            \$v3397\ := \$arr1452_ptr_take\;
            if \$v3397\(0) = '1' then
              \state\ <= q_wait3396;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3394;
            end if;
          when q_wait3400 =>
            \$v3401\ := \$arr1452_ptr_take\;
            if \$v3401\(0) = '1' then
              \state\ <= q_wait3400;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3398;
            end if;
          when q_wait3404 =>
            \$v3405\ := \$arr1451_ptr_take\;
            if \$v3405\(0) = '1' then
              \state\ <= q_wait3404;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1219\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1220\;
              \state\ <= pause_setI3402;
            end if;
          when q_wait3409 =>
            \$v3410\ := \$arr1451_ptr_take\;
            if \$v3410\(0) = '1' then
              \state\ <= q_wait3409;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1227\));
              \state\ <= pause_getI3407;
            end if;
          when q_wait3414 =>
            \$v3415\ := \$arr1452_ptr_take\;
            if \$v3415\(0) = '1' then
              \state\ <= q_wait3414;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3412;
            end if;
          when q_wait3418 =>
            \$v3419\ := \$arr1451_ptr_take\;
            if \$v3419\(0) = '1' then
              \state\ <= q_wait3418;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1233\));
              \state\ <= pause_getI3416;
            end if;
          when q_wait3423 =>
            \$v3424\ := \$arr1452_ptr_take\;
            if \$v3424\(0) = '1' then
              \state\ <= q_wait3423;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3421;
            end if;
          when q_wait3428 =>
            \$v3429\ := \$arr1452_ptr_take\;
            if \$v3429\(0) = '1' then
              \state\ <= q_wait3428;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3426;
            end if;
          when q_wait3436 =>
            \$v3437\ := \$arr1451_ptr_take\;
            if \$v3437\(0) = '1' then
              \state\ <= q_wait3436;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1255\));
              \state\ <= pause_getI3434;
            end if;
          when q_wait3441 =>
            \$v3442\ := \$arr1452_ptr_take\;
            if \$v3442\(0) = '1' then
              \state\ <= q_wait3441;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3439;
            end if;
          when q_wait3445 =>
            \$v3446\ := \$arr1451_ptr_take\;
            if \$v3446\(0) = '1' then
              \state\ <= q_wait3445;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1261\));
              \state\ <= pause_getI3443;
            end if;
          when q_wait3450 =>
            \$v3451\ := \$arr1452_ptr_take\;
            if \$v3451\(0) = '1' then
              \state\ <= q_wait3450;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3448;
            end if;
          when q_wait3454 =>
            \$v3455\ := \$arr1453_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 5;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v95\;
              \state\ <= pause_setI3452;
            end if;
          when q_wait3460 =>
            \$v3461\ := \$arr1452_ptr_take\;
            if \$v3461\(0) = '1' then
              \state\ <= q_wait3460;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3458;
            end if;
          when q_wait3464 =>
            \$v3465\ := \$arr1451_ptr_take\;
            if \$v3465\(0) = '1' then
              \state\ <= q_wait3464;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$74_result_after_f\;
              \state\ <= pause_setI3462;
            end if;
          when q_wait3470 =>
            \$v3471\ := \$arr1452_ptr_take\;
            if \$v3471\(0) = '1' then
              \state\ <= q_wait3470;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3468;
            end if;
          when q_wait3476 =>
            \$v3477\ := \$arr1451_ptr_take\;
            if \$v3477\(0) = '1' then
              \state\ <= q_wait3476;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3472\ := eclat_sub(\$1263_i\ & "00000000000000000000000000000001");
              \$v3473\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3472\ & "0010" & \$1263_i\ & "0001" & \$v3473\;
              \state\ <= pause_setI3474;
            end if;
          when q_wait3480 =>
            \$v3481\ := \$arr1451_ptr_take\;
            if \$v3481\(0) = '1' then
              \state\ <= q_wait3480;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1263_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$74_result_after_f\;
              \state\ <= pause_setI3478;
            end if;
          when q_wait3487 =>
            \$v3488\ := \$arr1452_ptr_take\;
            if \$v3488\(0) = '1' then
              \state\ <= q_wait3487;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3485;
            end if;
          when q_wait3505 =>
            \$v3506\ := \$arr1451_ptr_take\;
            if \$v3506\(0) = '1' then
              \state\ <= q_wait3505;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1300\));
              \state\ <= pause_getI3503;
            end if;
          when q_wait3510 =>
            \$v3511\ := \$arr1452_ptr_take\;
            if \$v3511\(0) = '1' then
              \state\ <= q_wait3510;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3508;
            end if;
          when q_wait3514 =>
            \$v3515\ := \$arr1452_ptr_take\;
            if \$v3515\(0) = '1' then
              \state\ <= q_wait3514;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3512;
            end if;
          when q_wait3518 =>
            \$v3519\ := \$arr1451_ptr_take\;
            if \$v3519\(0) = '1' then
              \state\ <= q_wait3518;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1272\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1273\;
              \state\ <= pause_setI3516;
            end if;
          when q_wait3523 =>
            \$v3524\ := \$arr1451_ptr_take\;
            if \$v3524\(0) = '1' then
              \state\ <= q_wait3523;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1280\));
              \state\ <= pause_getI3521;
            end if;
          when q_wait3528 =>
            \$v3529\ := \$arr1452_ptr_take\;
            if \$v3529\(0) = '1' then
              \state\ <= q_wait3528;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3526;
            end if;
          when q_wait3532 =>
            \$v3533\ := \$arr1451_ptr_take\;
            if \$v3533\(0) = '1' then
              \state\ <= q_wait3532;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1286\));
              \state\ <= pause_getI3530;
            end if;
          when q_wait3537 =>
            \$v3538\ := \$arr1452_ptr_take\;
            if \$v3538\(0) = '1' then
              \state\ <= q_wait3537;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3535;
            end if;
          when q_wait3542 =>
            \$v3543\ := \$arr1452_ptr_take\;
            if \$v3543\(0) = '1' then
              \state\ <= q_wait3542;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3540;
            end if;
          when q_wait3550 =>
            \$v3551\ := \$arr1451_ptr_take\;
            if \$v3551\(0) = '1' then
              \state\ <= q_wait3550;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1308\));
              \state\ <= pause_getI3548;
            end if;
          when q_wait3555 =>
            \$v3556\ := \$arr1452_ptr_take\;
            if \$v3556\(0) = '1' then
              \state\ <= q_wait3555;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3553;
            end if;
          when q_wait3559 =>
            \$v3560\ := \$arr1451_ptr_take\;
            if \$v3560\(0) = '1' then
              \state\ <= q_wait3559;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1314\));
              \state\ <= pause_getI3557;
            end if;
          when q_wait3564 =>
            \$v3565\ := \$arr1452_ptr_take\;
            if \$v3565\(0) = '1' then
              \state\ <= q_wait3564;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3562;
            end if;
          when q_wait3568 =>
            \$v3569\ := \$arr1453_ptr_take\;
            if \$v3569\(0) = '1' then
              \state\ <= q_wait3568;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 4;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v94\;
              \state\ <= pause_setI3566;
            end if;
          when q_wait3574 =>
            \$v3575\ := \$arr1452_ptr_take\;
            if \$v3575\(0) = '1' then
              \state\ <= q_wait3574;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3572;
            end if;
          when q_wait3579 =>
            \$v3580\ := \$arr1451_ptr_take\;
            if \$v3580\(0) = '1' then
              \state\ <= q_wait3579;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3576\ := "00000000000000000000000000000001";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3576\;
              \state\ <= pause_setI3577;
            end if;
          when q_wait3585 =>
            \$v3586\ := \$arr1452_ptr_take\;
            if \$v3586\(0) = '1' then
              \state\ <= q_wait3585;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3583;
            end if;
          when q_wait3591 =>
            \$v3592\ := \$arr1451_ptr_take\;
            if \$v3592\(0) = '1' then
              \state\ <= q_wait3591;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3587\ := eclat_sub(\$1316_i\ & "00000000000000000000000000000001");
              \$v3588\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3587\ & "0010" & \$1316_i\ & "0001" & \$v3588\;
              \state\ <= pause_setI3589;
            end if;
          when q_wait3596 =>
            \$v3597\ := \$arr1451_ptr_take\;
            if \$v3597\(0) = '1' then
              \state\ <= q_wait3596;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3593\ := "00000000000000000000000000000001";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1316_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$59_tos\(0 to 35) & \$61_y\ & "0001" & \$v3593\;
              \state\ <= pause_setI3594;
            end if;
          when q_wait3603 =>
            \$v3604\ := \$arr1452_ptr_take\;
            if \$v3604\(0) = '1' then
              \state\ <= q_wait3603;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3601;
            end if;
          when q_wait3607 =>
            \$v3608\ := \$arr1451_ptr_take\;
            if \$v3608\(0) = '1' then
              \state\ <= q_wait3607;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v79\));
              \state\ <= pause_getI3605;
            end if;
          when q_wait3612 =>
            \$v3613\ := \$arr1452_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3610;
            end if;
          when q_wait3617 =>
            \$v3618\ := \$arr1451_ptr_take\;
            if \$v3618\(0) = '1' then
              \state\ <= q_wait3617;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1333_i\));
              \state\ <= pause_getI3615;
            end if;
          when q_wait3628 =>
            \$v3629\ := \$arr1451_ptr_take\;
            if \$v3629\(0) = '1' then
              \state\ <= q_wait3628;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1367\));
              \state\ <= pause_getI3626;
            end if;
          when q_wait3633 =>
            \$v3634\ := \$arr1452_ptr_take\;
            if \$v3634\(0) = '1' then
              \state\ <= q_wait3633;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3631;
            end if;
          when q_wait3637 =>
            \$v3638\ := \$arr1452_ptr_take\;
            if \$v3638\(0) = '1' then
              \state\ <= q_wait3637;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3635;
            end if;
          when q_wait3641 =>
            \$v3642\ := \$arr1451_ptr_take\;
            if \$v3642\(0) = '1' then
              \state\ <= q_wait3641;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1339\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1340\;
              \state\ <= pause_setI3639;
            end if;
          when q_wait3646 =>
            \$v3647\ := \$arr1451_ptr_take\;
            if \$v3647\(0) = '1' then
              \state\ <= q_wait3646;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1347\));
              \state\ <= pause_getI3644;
            end if;
          when q_wait3651 =>
            \$v3652\ := \$arr1452_ptr_take\;
            if \$v3652\(0) = '1' then
              \state\ <= q_wait3651;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3649;
            end if;
          when q_wait3655 =>
            \$v3656\ := \$arr1451_ptr_take\;
            if \$v3656\(0) = '1' then
              \state\ <= q_wait3655;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1353\));
              \state\ <= pause_getI3653;
            end if;
          when q_wait3660 =>
            \$v3661\ := \$arr1452_ptr_take\;
            if \$v3661\(0) = '1' then
              \state\ <= q_wait3660;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3658;
            end if;
          when q_wait3665 =>
            \$v3666\ := \$arr1452_ptr_take\;
            if \$v3666\(0) = '1' then
              \state\ <= q_wait3665;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3663;
            end if;
          when q_wait3673 =>
            \$v3674\ := \$arr1451_ptr_take\;
            if \$v3674\(0) = '1' then
              \state\ <= q_wait3673;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1375\));
              \state\ <= pause_getI3671;
            end if;
          when q_wait3678 =>
            \$v3679\ := \$arr1452_ptr_take\;
            if \$v3679\(0) = '1' then
              \state\ <= q_wait3678;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3676;
            end if;
          when q_wait3682 =>
            \$v3683\ := \$arr1451_ptr_take\;
            if \$v3683\(0) = '1' then
              \state\ <= q_wait3682;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1381\));
              \state\ <= pause_getI3680;
            end if;
          when q_wait3687 =>
            \$v3688\ := \$arr1452_ptr_take\;
            if \$v3688\(0) = '1' then
              \state\ <= q_wait3687;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3685;
            end if;
          when q_wait3691 =>
            \$v3692\ := \$arr1453_ptr_take\;
            if \$v3692\(0) = '1' then
              \state\ <= q_wait3691;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 3;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v93\;
              \state\ <= pause_setI3689;
            end if;
          when q_wait3698 =>
            \$v3699\ := \$arr1452_ptr_take\;
            if \$v3699\(0) = '1' then
              \state\ <= q_wait3698;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3696;
            end if;
          when q_wait3702 =>
            \$v3703\ := \$arr1452_ptr_take\;
            if \$v3703\(0) = '1' then
              \state\ <= q_wait3702;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3700;
            end if;
          when q_wait3708 =>
            \$v3709\ := \$arr1451_ptr_take\;
            if \$v3709\(0) = '1' then
              \state\ <= q_wait3708;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3704\ := "00000000000000000000000000000000";
              \$v3705\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1383_x\ & "0001" & \$v3704\ & "0001" & \$v3705\;
              \state\ <= pause_setI3706;
            end if;
          when q_wait3714 =>
            \$v3715\ := \$arr1452_ptr_take\;
            if \$v3715\(0) = '1' then
              \state\ <= q_wait3714;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3712;
            end if;
          when q_wait3719 =>
            \$v3720\ := \$arr1451_ptr_take\;
            if \$v3720\(0) = '1' then
              \state\ <= q_wait3719;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3716\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1385_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1383_x\ & "0010" & \$1385_i\ & "0001" & \$v3716\;
              \state\ <= pause_setI3717;
            end if;
          when q_wait3726 =>
            \$v3727\ := \$arr1452_ptr_take\;
            if \$v3727\(0) = '1' then
              \state\ <= q_wait3726;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3724;
            end if;
          when q_wait3735 =>
            \$v3736\ := \$arr1451_ptr_take\;
            if \$v3736\(0) = '1' then
              \state\ <= q_wait3735;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1426\));
              \state\ <= pause_getI3733;
            end if;
          when q_wait3740 =>
            \$v3741\ := \$arr1452_ptr_take\;
            if \$v3741\(0) = '1' then
              \state\ <= q_wait3740;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3738;
            end if;
          when q_wait3744 =>
            \$v3745\ := \$arr1452_ptr_take\;
            if \$v3745\(0) = '1' then
              \state\ <= q_wait3744;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3742;
            end if;
          when q_wait3748 =>
            \$v3749\ := \$arr1451_ptr_take\;
            if \$v3749\(0) = '1' then
              \state\ <= q_wait3748;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1398\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1399\;
              \state\ <= pause_setI3746;
            end if;
          when q_wait3753 =>
            \$v3754\ := \$arr1451_ptr_take\;
            if \$v3754\(0) = '1' then
              \state\ <= q_wait3753;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1406\));
              \state\ <= pause_getI3751;
            end if;
          when q_wait3758 =>
            \$v3759\ := \$arr1452_ptr_take\;
            if \$v3759\(0) = '1' then
              \state\ <= q_wait3758;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3756;
            end if;
          when q_wait3762 =>
            \$v3763\ := \$arr1451_ptr_take\;
            if \$v3763\(0) = '1' then
              \state\ <= q_wait3762;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1412\));
              \state\ <= pause_getI3760;
            end if;
          when q_wait3767 =>
            \$v3768\ := \$arr1452_ptr_take\;
            if \$v3768\(0) = '1' then
              \state\ <= q_wait3767;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3765;
            end if;
          when q_wait3772 =>
            \$v3773\ := \$arr1452_ptr_take\;
            if \$v3773\(0) = '1' then
              \state\ <= q_wait3772;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3770;
            end if;
          when q_wait3780 =>
            \$v3781\ := \$arr1451_ptr_take\;
            if \$v3781\(0) = '1' then
              \state\ <= q_wait3780;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1434\));
              \state\ <= pause_getI3778;
            end if;
          when q_wait3785 =>
            \$v3786\ := \$arr1452_ptr_take\;
            if \$v3786\(0) = '1' then
              \state\ <= q_wait3785;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3783;
            end if;
          when q_wait3789 =>
            \$v3790\ := \$arr1451_ptr_take\;
            if \$v3790\(0) = '1' then
              \state\ <= q_wait3789;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1440\));
              \state\ <= pause_getI3787;
            end if;
          when q_wait3794 =>
            \$v3795\ := \$arr1452_ptr_take\;
            if \$v3795\(0) = '1' then
              \state\ <= q_wait3794;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3792;
            end if;
          when q_wait3803 =>
            \$v3804\ := \$arr1451_ptr_take\;
            if \$v3804\(0) = '1' then
              \state\ <= q_wait3803;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1472\));
              \state\ <= pause_getI3801;
            end if;
          when q_wait3808 =>
            \$v3809\ := \$arr1452_ptr_take\;
            if \$v3809\(0) = '1' then
              \state\ <= q_wait3808;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3806;
            end if;
          when q_wait3812 =>
            \$v3813\ := \$arr1452_ptr_take\;
            if \$v3813\(0) = '1' then
              \state\ <= q_wait3812;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3810;
            end if;
          when q_wait3816 =>
            \$v3817\ := \$arr1451_ptr_take\;
            if \$v3817\(0) = '1' then
              \state\ <= q_wait3816;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1444\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1445\;
              \state\ <= pause_setI3814;
            end if;
          when q_wait3821 =>
            \$v3822\ := \$arr1451_ptr_take\;
            if \$v3822\(0) = '1' then
              \state\ <= q_wait3821;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1452\));
              \state\ <= pause_getI3819;
            end if;
          when q_wait3826 =>
            \$v3827\ := \$arr1452_ptr_take\;
            if \$v3827\(0) = '1' then
              \state\ <= q_wait3826;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3824;
            end if;
          when q_wait3830 =>
            \$v3831\ := \$arr1451_ptr_take\;
            if \$v3831\(0) = '1' then
              \state\ <= q_wait3830;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1458\));
              \state\ <= pause_getI3828;
            end if;
          when q_wait3835 =>
            \$v3836\ := \$arr1452_ptr_take\;
            if \$v3836\(0) = '1' then
              \state\ <= q_wait3835;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3833;
            end if;
          when q_wait3840 =>
            \$v3841\ := \$arr1452_ptr_take\;
            if \$v3841\(0) = '1' then
              \state\ <= q_wait3840;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3838;
            end if;
          when q_wait3848 =>
            \$v3849\ := \$arr1451_ptr_take\;
            if \$v3849\(0) = '1' then
              \state\ <= q_wait3848;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1480\));
              \state\ <= pause_getI3846;
            end if;
          when q_wait3853 =>
            \$v3854\ := \$arr1452_ptr_take\;
            if \$v3854\(0) = '1' then
              \state\ <= q_wait3853;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3851;
            end if;
          when q_wait3857 =>
            \$v3858\ := \$arr1451_ptr_take\;
            if \$v3858\(0) = '1' then
              \state\ <= q_wait3857;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1486\));
              \state\ <= pause_getI3855;
            end if;
          when q_wait3862 =>
            \$v3863\ := \$arr1452_ptr_take\;
            if \$v3863\(0) = '1' then
              \state\ <= q_wait3862;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3860;
            end if;
          when q_wait3866 =>
            \$v3867\ := \$arr1453_ptr_take\;
            if \$v3867\(0) = '1' then
              \state\ <= q_wait3866;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 1;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v91\;
              \state\ <= pause_setI3864;
            end if;
          when q_wait3873 =>
            \$v3874\ := \$arr1452_ptr_take\;
            if \$v3874\(0) = '1' then
              \state\ <= q_wait3873;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3871;
            end if;
          when q_wait3877 =>
            \$v3878\ := \$arr1452_ptr_take\;
            if \$v3878\(0) = '1' then
              \state\ <= q_wait3877;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3875;
            end if;
          when q_wait3883 =>
            \$v3884\ := \$arr1451_ptr_take\;
            if \$v3884\(0) = '1' then
              \state\ <= q_wait3883;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3879\ := "00000000000000000000000000000000";
              \$v3880\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$76_result\ & "0001" & \$v3879\ & "0001" & \$v3880\;
              \state\ <= pause_setI3881;
            end if;
          when q_wait3889 =>
            \$v3890\ := \$arr1452_ptr_take\;
            if \$v3890\(0) = '1' then
              \state\ <= q_wait3889;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3887;
            end if;
          when q_wait3894 =>
            \$v3895\ := \$arr1451_ptr_take\;
            if \$v3895\(0) = '1' then
              \state\ <= q_wait3894;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3891\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1488_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$76_result\ & "0010" & \$1488_i\ & "0001" & \$v3891\;
              \state\ <= pause_setI3892;
            end if;
          when q_wait3901 =>
            \$v3902\ := \$arr1452_ptr_take\;
            if \$v3902\(0) = '1' then
              \state\ <= q_wait3901;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3899;
            end if;
          when q_wait3910 =>
            \$v3911\ := \$arr1451_ptr_take\;
            if \$v3911\(0) = '1' then
              \state\ <= q_wait3910;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1529\));
              \state\ <= pause_getI3908;
            end if;
          when q_wait3915 =>
            \$v3916\ := \$arr1452_ptr_take\;
            if \$v3916\(0) = '1' then
              \state\ <= q_wait3915;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3913;
            end if;
          when q_wait3919 =>
            \$v3920\ := \$arr1452_ptr_take\;
            if \$v3920\(0) = '1' then
              \state\ <= q_wait3919;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3917;
            end if;
          when q_wait3923 =>
            \$v3924\ := \$arr1451_ptr_take\;
            if \$v3924\(0) = '1' then
              \state\ <= q_wait3923;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1501\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1502\;
              \state\ <= pause_setI3921;
            end if;
          when q_wait3928 =>
            \$v3929\ := \$arr1451_ptr_take\;
            if \$v3929\(0) = '1' then
              \state\ <= q_wait3928;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1509\));
              \state\ <= pause_getI3926;
            end if;
          when q_wait3933 =>
            \$v3934\ := \$arr1452_ptr_take\;
            if \$v3934\(0) = '1' then
              \state\ <= q_wait3933;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3931;
            end if;
          when q_wait3937 =>
            \$v3938\ := \$arr1451_ptr_take\;
            if \$v3938\(0) = '1' then
              \state\ <= q_wait3937;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1515\));
              \state\ <= pause_getI3935;
            end if;
          when q_wait3942 =>
            \$v3943\ := \$arr1452_ptr_take\;
            if \$v3943\(0) = '1' then
              \state\ <= q_wait3942;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3940;
            end if;
          when q_wait3947 =>
            \$v3948\ := \$arr1452_ptr_take\;
            if \$v3948\(0) = '1' then
              \state\ <= q_wait3947;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3945;
            end if;
          when q_wait3955 =>
            \$v3956\ := \$arr1451_ptr_take\;
            if \$v3956\(0) = '1' then
              \state\ <= q_wait3955;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1537\));
              \state\ <= pause_getI3953;
            end if;
          when q_wait3960 =>
            \$v3961\ := \$arr1452_ptr_take\;
            if \$v3961\(0) = '1' then
              \state\ <= q_wait3960;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3958;
            end if;
          when q_wait3964 =>
            \$v3965\ := \$arr1451_ptr_take\;
            if \$v3965\(0) = '1' then
              \state\ <= q_wait3964;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1543\));
              \state\ <= pause_getI3962;
            end if;
          when q_wait3969 =>
            \$v3970\ := \$arr1452_ptr_take\;
            if \$v3970\(0) = '1' then
              \state\ <= q_wait3969;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3967;
            end if;
          when q_wait3973 =>
            \$v3974\ := \$arr1453_ptr_take\;
            if \$v3974\(0) = '1' then
              \state\ <= q_wait3973;
            else
              \$arr1453_ptr_take\(0) := '1';
              \$arr1453_ptr_write\ <= 0;
              \$arr1453_write_request\ <= '1';
              \$arr1453_write\ <= \$v89\;
              \state\ <= pause_setI3971;
            end if;
          when q_wait3979 =>
            \$v3980\ := \$arr1452_ptr_take\;
            if \$v3980\(0) = '1' then
              \state\ <= q_wait3979;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3977;
            end if;
          when q_wait3983 =>
            \$v3984\ := \$arr1451_ptr_take\;
            if \$v3984\(0) = '1' then
              \state\ <= q_wait3983;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
              \state\ <= pause_setI3981;
            end if;
          when q_wait3989 =>
            \$v3990\ := \$arr1452_ptr_take\;
            if \$v3990\(0) = '1' then
              \state\ <= q_wait3989;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI3987;
            end if;
          when q_wait3995 =>
            \$v3996\ := \$arr1451_ptr_take\;
            if \$v3996\(0) = '1' then
              \state\ <= q_wait3995;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$v3991\ := eclat_sub(\$1545_i\ & "00000000000000000000000000000001");
              \$v3992\ := "00000000000000000000000000000000";
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000010")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= "0010" & \$v3991\ & "0010" & \$1545_i\ & "0001" & \$v3992\;
              \state\ <= pause_setI3993;
            end if;
          when q_wait3999 =>
            \$v4000\ := \$arr1451_ptr_take\;
            if \$v4000\(0) = '1' then
              \state\ <= q_wait3999;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1545_i\ & "00000000000000000000000000000001")));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$67_z\ & \$66_y\ & \$65_x\;
              \state\ <= pause_setI3997;
            end if;
          when q_wait4006 =>
            \$v4007\ := \$arr1452_ptr_take\;
            if \$v4007\(0) = '1' then
              \state\ <= q_wait4006;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4004;
            end if;
          when q_wait4015 =>
            \$v4016\ := \$arr1451_ptr_take\;
            if \$v4016\(0) = '1' then
              \state\ <= q_wait4015;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1582\));
              \state\ <= pause_getI4013;
            end if;
          when q_wait4020 =>
            \$v4021\ := \$arr1452_ptr_take\;
            if \$v4021\(0) = '1' then
              \state\ <= q_wait4020;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4018;
            end if;
          when q_wait4024 =>
            \$v4025\ := \$arr1452_ptr_take\;
            if \$v4025\(0) = '1' then
              \state\ <= q_wait4024;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4022;
            end if;
          when q_wait4028 =>
            \$v4029\ := \$arr1451_ptr_take\;
            if \$v4029\(0) = '1' then
              \state\ <= q_wait4028;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1554\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1555\;
              \state\ <= pause_setI4026;
            end if;
          when q_wait4033 =>
            \$v4034\ := \$arr1451_ptr_take\;
            if \$v4034\(0) = '1' then
              \state\ <= q_wait4033;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1562\));
              \state\ <= pause_getI4031;
            end if;
          when q_wait4038 =>
            \$v4039\ := \$arr1452_ptr_take\;
            if \$v4039\(0) = '1' then
              \state\ <= q_wait4038;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4036;
            end if;
          when q_wait4042 =>
            \$v4043\ := \$arr1451_ptr_take\;
            if \$v4043\(0) = '1' then
              \state\ <= q_wait4042;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1568\));
              \state\ <= pause_getI4040;
            end if;
          when q_wait4047 =>
            \$v4048\ := \$arr1452_ptr_take\;
            if \$v4048\(0) = '1' then
              \state\ <= q_wait4047;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4045;
            end if;
          when q_wait4052 =>
            \$v4053\ := \$arr1452_ptr_take\;
            if \$v4053\(0) = '1' then
              \state\ <= q_wait4052;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4050;
            end if;
          when q_wait4060 =>
            \$v4061\ := \$arr1451_ptr_take\;
            if \$v4061\(0) = '1' then
              \state\ <= q_wait4060;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1590\));
              \state\ <= pause_getI4058;
            end if;
          when q_wait4065 =>
            \$v4066\ := \$arr1452_ptr_take\;
            if \$v4066\(0) = '1' then
              \state\ <= q_wait4065;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4063;
            end if;
          when q_wait4069 =>
            \$v4070\ := \$arr1451_ptr_take\;
            if \$v4070\(0) = '1' then
              \state\ <= q_wait4069;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1596\));
              \state\ <= pause_getI4067;
            end if;
          when q_wait4074 =>
            \$v4075\ := \$arr1452_ptr_take\;
            if \$v4075\(0) = '1' then
              \state\ <= q_wait4074;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4072;
            end if;
          when q_wait4083 =>
            \$v4084\ := \$arr1451_ptr_take\;
            if \$v4084\(0) = '1' then
              \state\ <= q_wait4083;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1628\));
              \state\ <= pause_getI4081;
            end if;
          when q_wait4088 =>
            \$v4089\ := \$arr1452_ptr_take\;
            if \$v4089\(0) = '1' then
              \state\ <= q_wait4088;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4086;
            end if;
          when q_wait4092 =>
            \$v4093\ := \$arr1452_ptr_take\;
            if \$v4093\(0) = '1' then
              \state\ <= q_wait4092;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4090;
            end if;
          when q_wait4096 =>
            \$v4097\ := \$arr1451_ptr_take\;
            if \$v4097\(0) = '1' then
              \state\ <= q_wait4096;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1600\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1601\;
              \state\ <= pause_setI4094;
            end if;
          when q_wait4101 =>
            \$v4102\ := \$arr1451_ptr_take\;
            if \$v4102\(0) = '1' then
              \state\ <= q_wait4101;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1608\));
              \state\ <= pause_getI4099;
            end if;
          when q_wait4106 =>
            \$v4107\ := \$arr1452_ptr_take\;
            if \$v4107\(0) = '1' then
              \state\ <= q_wait4106;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4104;
            end if;
          when q_wait4110 =>
            \$v4111\ := \$arr1451_ptr_take\;
            if \$v4111\(0) = '1' then
              \state\ <= q_wait4110;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1614\));
              \state\ <= pause_getI4108;
            end if;
          when q_wait4115 =>
            \$v4116\ := \$arr1452_ptr_take\;
            if \$v4116\(0) = '1' then
              \state\ <= q_wait4115;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4113;
            end if;
          when q_wait4120 =>
            \$v4121\ := \$arr1452_ptr_take\;
            if \$v4121\(0) = '1' then
              \state\ <= q_wait4120;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4118;
            end if;
          when q_wait4128 =>
            \$v4129\ := \$arr1451_ptr_take\;
            if \$v4129\(0) = '1' then
              \state\ <= q_wait4128;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1636\));
              \state\ <= pause_getI4126;
            end if;
          when q_wait4133 =>
            \$v4134\ := \$arr1452_ptr_take\;
            if \$v4134\(0) = '1' then
              \state\ <= q_wait4133;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4131;
            end if;
          when q_wait4137 =>
            \$v4138\ := \$arr1451_ptr_take\;
            if \$v4138\(0) = '1' then
              \state\ <= q_wait4137;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1642\));
              \state\ <= pause_getI4135;
            end if;
          when q_wait4142 =>
            \$v4143\ := \$arr1452_ptr_take\;
            if \$v4143\(0) = '1' then
              \state\ <= q_wait4142;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4140;
            end if;
          when q_wait4151 =>
            \$v4152\ := \$arr1451_ptr_take\;
            if \$v4152\(0) = '1' then
              \state\ <= q_wait4151;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1674\));
              \state\ <= pause_getI4149;
            end if;
          when q_wait4156 =>
            \$v4157\ := \$arr1452_ptr_take\;
            if \$v4157\(0) = '1' then
              \state\ <= q_wait4156;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4154;
            end if;
          when q_wait4160 =>
            \$v4161\ := \$arr1452_ptr_take\;
            if \$v4161\(0) = '1' then
              \state\ <= q_wait4160;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4158;
            end if;
          when q_wait4164 =>
            \$v4165\ := \$arr1451_ptr_take\;
            if \$v4165\(0) = '1' then
              \state\ <= q_wait4164;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr_write\ <= to_integer(unsigned(\$1646\));
              \$arr1451_write_request\ <= '1';
              \$arr1451_write\ <= \$1647\;
              \state\ <= pause_setI4162;
            end if;
          when q_wait4169 =>
            \$v4170\ := \$arr1451_ptr_take\;
            if \$v4170\(0) = '1' then
              \state\ <= q_wait4169;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1654\));
              \state\ <= pause_getI4167;
            end if;
          when q_wait4174 =>
            \$v4175\ := \$arr1452_ptr_take\;
            if \$v4175\(0) = '1' then
              \state\ <= q_wait4174;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4172;
            end if;
          when q_wait4178 =>
            \$v4179\ := \$arr1451_ptr_take\;
            if \$v4179\(0) = '1' then
              \state\ <= q_wait4178;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1660\));
              \state\ <= pause_getI4176;
            end if;
          when q_wait4183 =>
            \$v4184\ := \$arr1452_ptr_take\;
            if \$v4184\(0) = '1' then
              \state\ <= q_wait4183;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4181;
            end if;
          when q_wait4188 =>
            \$v4189\ := \$arr1452_ptr_take\;
            if \$v4189\(0) = '1' then
              \state\ <= q_wait4188;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4186;
            end if;
          when q_wait4196 =>
            \$v4197\ := \$arr1451_ptr_take\;
            if \$v4197\(0) = '1' then
              \state\ <= q_wait4196;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1682\));
              \state\ <= pause_getI4194;
            end if;
          when q_wait4201 =>
            \$v4202\ := \$arr1452_ptr_take\;
            if \$v4202\(0) = '1' then
              \state\ <= q_wait4201;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4199;
            end if;
          when q_wait4205 =>
            \$v4206\ := \$arr1451_ptr_take\;
            if \$v4206\(0) = '1' then
              \state\ <= q_wait4205;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$1688\));
              \state\ <= pause_getI4203;
            end if;
          when q_wait4210 =>
            \$v4211\ := \$arr1452_ptr_take\;
            if \$v4211\(0) = '1' then
              \state\ <= q_wait4210;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4208;
            end if;
          when q_wait4214 =>
            \$v4215\ := \$arr1451_ptr_take\;
            if \$v4215\(0) = '1' then
              \state\ <= q_wait4214;
            else
              \$arr1451_ptr_take\(0) := '1';
              \$arr1451_ptr\ <= to_integer(unsigned(\$v17\));
              \state\ <= pause_getI4212;
            end if;
          when q_wait4219 =>
            \$v4220\ := \$arr1452_ptr_take\;
            if \$v4220\(0) = '1' then
              \state\ <= q_wait4219;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr\ <= 1;
              \state\ <= pause_getI4217;
            end if;
          when q_wait4223 =>
            \$v4224\ := \$arr1452_ptr_take\;
            if \$v4224\(0) = '1' then
              \state\ <= q_wait4223;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 4;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= pos;
              \state\ <= pause_setI4221;
            end if;
          when q_wait4227 =>
            \$v4228\ := \$arr1452_ptr_take\;
            if \$v4228\(0) = '1' then
              \state\ <= q_wait4227;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 3;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= stbl;
              \state\ <= pause_setI4225;
            end if;
          when q_wait4231 =>
            \$v4232\ := \$arr1452_ptr_take\;
            if \$v4232\(0) = '1' then
              \state\ <= q_wait4231;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 2;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= st;
              \state\ <= pause_setI4229;
            end if;
          when q_wait4235 =>
            \$v4236\ := \$arr1452_ptr_take\;
            if \$v4236\(0) = '1' then
              \state\ <= q_wait4235;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 1;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= sp;
              \state\ <= pause_setI4233;
            end if;
          when q_wait4239 =>
            \$v4240\ := \$arr1452_ptr_take\;
            if \$v4240\(0) = '1' then
              \state\ <= q_wait4239;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 0;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= pc;
              \state\ <= pause_setI4237;
            end if;
          when compute1456 =>
            rdy1455 := eclat_false;
            pc := eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
            sp := X"000" & X"15f90";
            st := eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
            stbl := eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
            pos := "00000000000000000000000000000000";
            \$v4240\ := \$arr1452_ptr_take\;
            if \$v4240\(0) = '1' then
              \state\ <= q_wait4239;
            else
              \$arr1452_ptr_take\(0) := '1';
              \$arr1452_ptr_write\ <= 0;
              \$arr1452_write_request\ <= '1';
              \$arr1452_write\ <= pc;
              \state\ <= pause_setI4237;
            end if;
          end case;
          
          result <= result1454;
          rdy <= rdy1455;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
