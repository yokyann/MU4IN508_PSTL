-- code generated from the following source code:
--   ../RibbitVm/fail.ecl
--   ../RibbitVm/vm.ecl
--
-- with the following command:
--
--    ./eclat ../RibbitVm/fail.ecl ../RibbitVm/vm.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute3408, \$1069_list_tail637\, \$1070_get_int640\, \$1072_rest_loop668\, \$1073_loop667\, \$1113_forever6893378\, \$1122_forever6893379\, \$1134_forever6893380\, \$1143_forever6893381\, \$1152_forever6893382\, \$1169_forever6893383\, \$1178_forever6893384\, \$1190_forever6893385\, \$1199_forever6893386\, \$1208_forever6893387\, \$1225_forever6893388\, \$1234_forever6893389\, \$1246_forever6893390\, \$1255_forever6893391\, \$1264_forever6893392\, \$1281_forever6893393\, \$1290_forever6893394\, \$1302_forever6893395\, \$1311_forever6893396\, \$1320_forever6893397\, \$1371_show_rib6323365\, \$1388_forever6893337\, \$1400_forever6893366\, \$1410_forever6893367\, \$1418_forever6893368\, \$1423_print_value6133369\, \$1433_forever6893370\, \$1450_forever6893371\, \$1458_forever6893372\, \$1464_loop6693373\, \$1473_forever6893356\, \$1481_forever6893360\, \$1515_forever6893374\, \$1525_forever6893375\, \$1534_forever6893376\, \$1546_forever6893377\, \$1599_forever6893361\, \$1609_forever6893362\, \$1618_forever6893363\, \$1630_forever6893364\, \$1669_forever6893338\, \$1684_forever6893339\, \$373_forever6893335\, \$373_forever6893336\, \$373_forever6893337\, \$373_forever6893358\, \$411_show_rib6323357\, \$411_show_rib6323359\, pause_getI3413, pause_getI3421, pause_getI3431, pause_getI3435, pause_getI3439, pause_getI3443, pause_getI3456, pause_getI3468, pause_getI3474, pause_getI3483, pause_getI3489, pause_getI3493, pause_getI3497, pause_getI3512, pause_getI3524, pause_getI3529, pause_getI3534, pause_getI3547, pause_getI3559, pause_getI3565, pause_getI3574, pause_getI3580, pause_getI3584, pause_getI3588, pause_getI3601, pause_getI3610, pause_getI3629, pause_getI3637, pause_getI3646, pause_getI3656, pause_getI3660, pause_getI3669, pause_getI3676, pause_getI3682, pause_getI3696, pause_getI3706, pause_getI3721, pause_getI3733, pause_getI3739, pause_getI3756, pause_getI3762, pause_getI3774, pause_getI3782, pause_getI3788, pause_getI3800, pause_getI3806, pause_getI3818, pause_getI3826, pause_getI3832, pause_getI3844, pause_getI3850, pause_getI3862, pause_getI3870, pause_getI3876, pause_getI3888, pause_getI3894, pause_getI3906, pause_getI3914, pause_getI3920, pause_getI3928, pause_getI3936, pause_getI3946, pause_getI3954, pause_getII3414, pause_getII3422, pause_getII3432, pause_getII3436, pause_getII3440, pause_getII3444, pause_getII3457, pause_getII3469, pause_getII3475, pause_getII3484, pause_getII3490, pause_getII3494, pause_getII3498, pause_getII3513, pause_getII3525, pause_getII3530, pause_getII3535, pause_getII3548, pause_getII3560, pause_getII3566, pause_getII3575, pause_getII3581, pause_getII3585, pause_getII3589, pause_getII3602, pause_getII3611, pause_getII3630, pause_getII3638, pause_getII3647, pause_getII3657, pause_getII3661, pause_getII3670, pause_getII3677, pause_getII3683, pause_getII3697, pause_getII3707, pause_getII3722, pause_getII3734, pause_getII3740, pause_getII3757, pause_getII3763, pause_getII3775, pause_getII3783, pause_getII3789, pause_getII3801, pause_getII3807, pause_getII3819, pause_getII3827, pause_getII3833, pause_getII3845, pause_getII3851, pause_getII3863, pause_getII3871, pause_getII3877, pause_getII3889, pause_getII3895, pause_getII3907, pause_getII3915, pause_getII3921, pause_getII3929, pause_getII3937, pause_getII3947, pause_getII3955, pause_setI3427, pause_setI3447, pause_setI3452, pause_setI3460, pause_setI3504, pause_setI3508, pause_setI3516, pause_setI3520, pause_setI3538, pause_setI3543, pause_setI3551, pause_setI3614, pause_setI3621, pause_setI3652, pause_setI3664, pause_setI3748, pause_setI3767, pause_setI3792, pause_setI3811, pause_setI3836, pause_setI3855, pause_setI3880, pause_setI3899, pause_setI3924, pause_setI3932, pause_setI3940, pause_setI3950, pause_setI3958, pause_setI3965, pause_setI3972, pause_setI3979, pause_setI3986, pause_setI3990, pause_setI3994, pause_setI3998, pause_setI4002, pause_setI4006, pause_setI4010, pause_setI4014, pause_setI4018, pause_setI4022, pause_setI4026, pause_setI4030, pause_setII3428, pause_setII3448, pause_setII3453, pause_setII3461, pause_setII3505, pause_setII3509, pause_setII3517, pause_setII3521, pause_setII3539, pause_setII3544, pause_setII3552, pause_setII3615, pause_setII3622, pause_setII3653, pause_setII3665, pause_setII3749, pause_setII3768, pause_setII3793, pause_setII3812, pause_setII3837, pause_setII3856, pause_setII3881, pause_setII3900, pause_setII3925, pause_setII3933, pause_setII3941, pause_setII3951, pause_setII3959, pause_setII3966, pause_setII3973, pause_setII3980, pause_setII3987, pause_setII3991, pause_setII3995, pause_setII3999, pause_setII4003, pause_setII4007, pause_setII4011, pause_setII4015, pause_setII4019, pause_setII4023, pause_setII4027, pause_setII4031, q_wait3415, q_wait3423, q_wait3429, q_wait3433, q_wait3437, q_wait3441, q_wait3445, q_wait3449, q_wait3454, q_wait3458, q_wait3462, q_wait3470, q_wait3476, q_wait3485, q_wait3491, q_wait3495, q_wait3499, q_wait3506, q_wait3510, q_wait3514, q_wait3518, q_wait3522, q_wait3526, q_wait3531, q_wait3536, q_wait3540, q_wait3545, q_wait3549, q_wait3553, q_wait3561, q_wait3567, q_wait3576, q_wait3582, q_wait3586, q_wait3590, q_wait3603, q_wait3612, q_wait3616, q_wait3623, q_wait3631, q_wait3639, q_wait3648, q_wait3654, q_wait3658, q_wait3662, q_wait3666, q_wait3671, q_wait3678, q_wait3684, q_wait3698, q_wait3708, q_wait3723, q_wait3735, q_wait3741, q_wait3750, q_wait3758, q_wait3764, q_wait3769, q_wait3776, q_wait3784, q_wait3790, q_wait3794, q_wait3802, q_wait3808, q_wait3813, q_wait3820, q_wait3828, q_wait3834, q_wait3838, q_wait3846, q_wait3852, q_wait3857, q_wait3864, q_wait3872, q_wait3878, q_wait3882, q_wait3890, q_wait3896, q_wait3901, q_wait3908, q_wait3916, q_wait3922, q_wait3926, q_wait3930, q_wait3934, q_wait3938, q_wait3942, q_wait3948, q_wait3952, q_wait3956, q_wait3960, q_wait3967, q_wait3974, q_wait3981, q_wait3988, q_wait3992, q_wait3996, q_wait4000, q_wait4004, q_wait4008, q_wait4012, q_wait4016, q_wait4020, q_wait4024, q_wait4028, q_wait4032);
  signal \state\: t_state;
  type array_value_32 is array (natural range <>) of value(0 to 31);
  type array_value_108 is array (natural range <>) of value(0 to 107);
  signal arr3398 : array_value_32(0 to 8999) := (others => (others => '0'));
  signal \$arr3398_value\ : value(0 to 31);
  signal \$arr3398_ptr\ : natural range 0 to 8999;
  signal \$arr3398_ptr_write\ : natural range 0 to 8999;
  signal \$arr3398_write\ : value(0 to 31);
  signal \$arr3398_write_request\ : std_logic := '0';
  signal arr3399 : array_value_108(0 to 8999) := (others => (others => '0'));
  signal \$arr3399_value\ : value(0 to 107);
  signal \$arr3399_ptr\ : natural range 0 to 8999;
  signal \$arr3399_ptr_write\ : natural range 0 to 8999;
  signal \$arr3399_write\ : value(0 to 107);
  signal \$arr3399_write_request\ : std_logic := '0';
  signal arr3400 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3400_value\ : value(0 to 31);
  signal \$arr3400_ptr\ : natural range 0 to 0;
  signal \$arr3400_ptr_write\ : natural range 0 to 0;
  signal \$arr3400_write\ : value(0 to 31);
  signal \$arr3400_write_request\ : std_logic := '0';
  signal arr3401 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3401_value\ : value(0 to 31);
  signal \$arr3401_ptr\ : natural range 0 to 0;
  signal \$arr3401_ptr_write\ : natural range 0 to 0;
  signal \$arr3401_write\ : value(0 to 31);
  signal \$arr3401_write_request\ : std_logic := '0';
  signal arr3402 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3402_value\ : value(0 to 31);
  signal \$arr3402_ptr\ : natural range 0 to 0;
  signal \$arr3402_ptr_write\ : natural range 0 to 0;
  signal \$arr3402_write\ : value(0 to 31);
  signal \$arr3402_write_request\ : std_logic := '0';
  signal arr3403 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3403_value\ : value(0 to 31);
  signal \$arr3403_ptr\ : natural range 0 to 0;
  signal \$arr3403_ptr_write\ : natural range 0 to 0;
  signal \$arr3403_write\ : value(0 to 31);
  signal \$arr3403_write_request\ : std_logic := '0';
  signal arr3404 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3404_value\ : value(0 to 31);
  signal \$arr3404_ptr\ : natural range 0 to 0;
  signal \$arr3404_ptr_write\ : natural range 0 to 0;
  signal \$arr3404_write\ : value(0 to 31);
  signal \$arr3404_write_request\ : std_logic := '0';
  signal arr3405 : array_value_32(0 to 5) := (others => (others => '0'));
  signal \$arr3405_value\ : value(0 to 31);
  signal \$arr3405_ptr\ : natural range 0 to 5;
  signal \$arr3405_ptr_write\ : natural range 0 to 5;
  signal \$arr3405_write\ : value(0 to 31);
  signal \$arr3405_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3398_write_request\ = '1' then
                    arr3398(\$arr3398_ptr_write\) <= \$arr3398_write\;
                  else
                   \$arr3398_value\ <= arr3398(\$arr3398_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3399_write_request\ = '1' then
                    arr3399(\$arr3399_ptr_write\) <= \$arr3399_write\;
                  else
                   \$arr3399_value\ <= arr3399(\$arr3399_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3400_write_request\ = '1' then
                    arr3400(\$arr3400_ptr_write\) <= \$arr3400_write\;
                  else
                   \$arr3400_value\ <= arr3400(\$arr3400_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3401_write_request\ = '1' then
                    arr3401(\$arr3401_ptr_write\) <= \$arr3401_write\;
                  else
                   \$arr3401_value\ <= arr3401(\$arr3401_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3402_write_request\ = '1' then
                    arr3402(\$arr3402_ptr_write\) <= \$arr3402_write\;
                  else
                   \$arr3402_value\ <= arr3402(\$arr3402_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3403_write_request\ = '1' then
                    arr3403(\$arr3403_ptr_write\) <= \$arr3403_write\;
                  else
                   \$arr3403_value\ <= arr3403(\$arr3403_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3404_write_request\ = '1' then
                    arr3404(\$arr3404_ptr_write\) <= \$arr3404_write\;
                  else
                   \$arr3404_value\ <= arr3404(\$arr3404_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3405_write_request\ = '1' then
                    arr3405(\$arr3405_ptr_write\) <= \$arr3405_write\;
                  else
                   \$arr3405_value\ <= arr3405(\$arr3405_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$v3480\, \$v3867\, \$1575\, \$1229\, \$v3717\, \$1213_car\, 
               \$1501\, \$v3641\, \$v3823\, \$1688\, \$v3797\, \$v3786\, 
               \$1467_tag\, \$1463\, \$1520\, \$v3816\, \$v3904\, \$v3626\, 
               \$v3737\, \$1438_k\, \$v3713\, \$v402\, \$1276\, \$1393\, 
               \$1333\, \$v3727\, \$v3563\, \$v3841\, \$v3760\, \$v3892\, 
               \$v3772\, \$v3633\, \$1585\, \$v3556\, \$1157_car\, \$v3465\, 
               \$1491\, \$v3710\, \$1444\, \$v3619\, \$v3848\, \$v3411\, 
               \$1604\, \$1269_car\, \$v3680\, \$1422\, \$v3918\, \$1445\, 
               \$1147\, \$v3885\, \$1117\, \$v3593\, \$1539\, \$v3578\, 
               \$1259\, \$1101_car\, \$v3725\, \$v3673\, \$v3650\, \$v3860\, 
               \$v3911\, \$v3597\, \$v3692\, \$v3419\, \$1108\, \$v3745\, 
               \$v3830\, \$v3730\, \$v3700\, \$1464_loop6693373_result\, 
               \$1541\, \$v3804\, \$1464_loop6693373_arg\, \$1285\, \$1625\, 
               \$v3605\, \$v3702\, \$1529\, \$1623\, \$1164\, 
               \$1423_print_value6133369_arg\, \$v3874\, \$v3607\, \$v3643\, 
               \$v3688\, \$v3472\, \$1315\, \$1203\, \$1220\, \$v3571\, 
               \$1613\, \$1173\, \$v3753\, \$1405\, \$v3779\, \$v3487\ : value(0 to 35) := (others => '0');
      variable \$1650\, \$1677\, \$1656\, \$1069_list_tail637_arg\ : value(0 to 63) := (others => '0');
      variable \$1072_rest_loop668_arg\ : value(0 to 131) := (others => '0');
      variable \$v3420\, \$v3773\, \$v3886\, \$v3893\, \$v3651\, \$v3738\, 
               \$v3693\, \$v3606\, \$v3849\, \$v3674\, \$v3473\, \$v3642\, 
               \$v3761\, \$v3466\, \$v3868\, \$v3805\, \$v3817\, \$v3634\, 
               \$v3481\, \$v3557\, \$v3728\, \$v3579\, \$v3701\, \$v3689\, 
               \$v3831\, \$v3488\, \$v3620\, \$v3905\, \$v3572\, \$v3726\, 
               \$v3875\, \$v3731\, \$v3711\, \$v3919\, \$v3644\, \$v3564\, 
               \$v3681\, \$v3798\, \$v3594\, \$v3608\, \$v3787\, \$v3780\, 
               \$v3824\, \$v3754\, \$v3412\, \$v3598\, \$v3714\, \$v3627\, 
               \$v3746\, \$v3718\, \$v3861\, \$v3842\, \$v3912\, \$v3703\ : value(0 to 3) := (others => '0');
      variable \$v4017\, \$v3569\, \$v3507\, \$v3426\, \$v3532\, \$v3715\, 
               \$v3417\, \$v3424\, \$v3736\, \$v3609\, \$v4013\, \$1665\, 
               \$v3814\, \$v3416\, \$v3463\, \$v3923\, \$v3679\, 
               \$1423_print_value6133369_result\, \$v3927\, \$v3821\, 
               \$v3477\, \$1371_show_rib6323365_result\, \$v3989\, \$v3729\, 
               \$v3471\, \$v3568\, \$v3803\, \$v3770\, \$v3550\, \$v3742\, 
               \$v3902\, \$v3617\, \$v3724\, \$v3595\, \$v3519\, \$v3865\, 
               \$1595\, \$v3982\, \$v3511\, \$v3546\, \$v3785\, \$v3809\, 
               \$v3939\, \$v3537\, \$v3649\, \$v3829\, \$v3604\, \$v3968\, 
               \$v3909\, \$v3791\, \$913\, \$v3917\, \$v3957\, \$v3751\, 
               \$v3847\, \$v3975\, \$v3879\, \$v3425\, \$v3897\, \$v3672\, 
               \$v3663\, \$v3765\, \$v3478\, \$v4021\, \$v3699\, \$v3777\, 
               \$v3583\, \$v3997\, rdy3407, \$v3655\, \$v3577\, \$v4005\, 
               \$v3935\, \$v3515\, \$v3533\, \$v3554\, \$v3858\, \$v3931\, 
               \$v3961\, \$v4029\, \$v3492\, \$v4001\, \$v3430\, \$v4033\, 
               \$v3759\, \$v3704\, result3406, \$1382\, \$v3591\, \$v3747\, 
               \$411_show_rib6323357_result\, \$1511\, \$v3835\, \$v3839\, 
               \$v3486\, \$v3496\, \$v3459\, \$v3943\, \$v3853\, \$v3442\, 
               \$v3690\, \$411_show_rib6323359_result\, \$v3949\, \$v4009\, 
               \$v3873\, \$v3709\, \$v4025\, \$v3434\, \$v3500\, \$v3659\, 
               \$v3523\, \$v3640\, \$v3953\, \$v3883\, \$v3667\, \$v3450\, 
               \$v3527\, \$v3541\, \$v3743\, \$v3455\, \$v3446\, \$v3562\, 
               \$v3891\, \$v3632\, \$v3993\, \$v3624\, \$v3685\, \$1437\, 
               \$v3795\, \$v3438\, \$v3587\, \$v3613\ : value(0 to 0) := (others => '0');
      variable \$1073_loop667_arg\ : value(0 to 171) := (others => '0');
      variable \$1690\, \$v1685\, \$1570\, \$1486\, \$v1675\, \$1439\, 
               \$v3315\, \$v2920\, \$v1723\, \$v3302\, \$v2950\, \$1214\, 
               \$1494\, \$1328\, \$v1713\, \$1270\, \$1490\, \$v1704\, 
               \$v2976\, \$v2929\, \$v2985\, \$v2925\, \$1673\, \$1102\, 
               \$1443\, \$1158\, \$v1666\, \$v1694\, \$v2916\, \$v2972\, 
               \$1327\, \$v2989\, \$1578\, \$v1656\, \$v2946\ : value(0 to 107) := (others => '0');
      variable \$411_show_rib6323357_arg\, \$1371_show_rib6323365_arg\, 
               \$411_show_rib6323359_arg\, \$1370\ : value(0 to 99) := (others => '0');
      variable \$1295\, \$1634\, \$v3962\, \$v3778\, \$1404\, \$v3635\, 
               \$v3687\, \$1238\, \$v3945\, \$v3744\, \$v3479\, \$v3903\, 
               \$1614_t\, \$1275\, \$v3502\, \$1648_x\, \$v3599\, \$1569\, 
               \$v3694\, \$1551\, \$1394\, \$1212\, \$1182\, \$1126\, 
               \$v3815\, \$1239\, \$1148_t\, \$v3636\, \$v3695\, \$1118_t\, 
               \$v3810\, \$1395\, \$1542_t\, \$1429_t\, \$v3971\, \$v3592\, 
               \$1251_i\, \$v3796\, \$v3720\, \$1306\, \$v3732\, \$1163\, 
               \$1138\, \$v3859\, \$1587\, \$v3977\, \$1530_t\, \$1538\, 
               \$v3501\, \$v3503\, \$v3558\, \$1588_i\, \$v3528\, \$1622\, 
               \$1428_i\, \$1657\, \$1396_i\, \$v3410\, \$v3970\, \$v3625\, 
               \$v3910\, \$v3409\, \$v3884\, \$v3766\, \$1550\, \$1414_t\, 
               \$1477_t\, \$1230_t\, \$1605_i\, \$v3840\, \$v3887\, \$v3573\, 
               \$914\, \$1316_t\, \$1130_i\, \$1156\, \$v3570\, \$1485\, 
               \$v3596\, \$1454_t\, \$v3716\, \$1655\, \$v3755\, \$v3822\, 
               \$1492\, \$1653_c\, \$1658\, \$v3825\, \$v3467\, \$v3618\, 
               \$1049_i\, \$v3691\, \$1139_i\, \$v3675\, \$1260_t\, \$v3976\, 
               \$1384_i\, \$v3628\, \$1165_i\, \$1183\, 
               \$1070_get_int640_arg\, \$v3668\, \$1107\, \$v3854\, 
               \$1571_i\, \$v3983\, \$1127\, \$v3984\, \$1651\, \$1277_i\, 
               \$v3869\, \$v3719\, \$v3418\, \$v3542\, \$v3964\, \$v3771\, 
               \$v3799\, \$1009_t\, \$1680_i\, \$1577\, \$1109_i\, \$v3985\, 
               \$1053_i\, \$v3645\, \$1242_i\, \$v3712\, \$v3482\, \$1325\, 
               \$1383\, \$1204_t\, \$1519\, \$v3464\, \$v3781\, \$1186_i\, 
               \$v3866\, \$v3944\, \$1504_i\, \$1446_t\, \$1194\, \$v3963\, 
               \$1336\, \$1521_i\, \$1503\, \$v3705\, \$1250\, \$v3752\, 
               \$v3978\, \$1603\, \$1294\, \$v3898\, \$1678\, \$1426_t\, 
               \$1307_i\, \$911_i\, \$1298_i\, \$1638_x\, \$v3843\, 
               \$1626_t\, \$1268\, \$1174_t\, \$1380_i\, \$1324\, \$1286_t\, 
               \$v3600\, \$v3451\, \$v3686\, \$1326\, \$1219\, \$1406_i\, 
               \$v3969\, \$1195_i\, \$1337\, \$1221_i\, \$1635\, \$v3913\, 
               \$v3555\ : value(0 to 31) := (others => '0');
      variable \$1584\, \$1500\ : value(0 to 67) := (others => '0');
      variable \$arr3398_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3399_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3400_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3401_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3402_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3403_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3404_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3405_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v3555\); default_zero(\$v3613\); 
          default_zero(\$1370\); default_zero(\$v3587\); 
          default_zero(\$v3913\); default_zero(\$1635\); 
          default_zero(\$v3438\); default_zero(\$1221_i\); 
          default_zero(\$v3487\); default_zero(\$v3795\); 
          default_zero(\$1337\); default_zero(\$1437\); 
          default_zero(\$v3779\); default_zero(\$v2946\); 
          default_zero(\$v3703\); default_zero(\$v3912\); 
          default_zero(\$1195_i\); default_zero(\$v3685\); 
          default_zero(\$v3969\); default_zero(\$v3624\); 
          default_zero(\$1069_list_tail637_arg\); default_zero(\$1405\); 
          default_zero(\$v3753\); default_zero(\$v3993\); 
          default_zero(\$v3632\); default_zero(\$v3842\); 
          default_zero(\$1406_i\); default_zero(\$1219\); 
          default_zero(\$1173\); default_zero(\$v1656\); 
          default_zero(\$1326\); default_zero(\$v3686\); 
          default_zero(\$1613\); default_zero(\$v3451\); 
          default_zero(\$v3600\); default_zero(\$v3861\); 
          default_zero(\$1578\); default_zero(\$v3891\); 
          default_zero(\$1286_t\); default_zero(\$1324\); 
          default_zero(\$v3571\); default_zero(\$v3562\); 
          default_zero(\$1380_i\); default_zero(\$1174_t\); 
          default_zero(\$v3446\); default_zero(\$1268\); 
          default_zero(\$v3455\); default_zero(\$v3718\); 
          default_zero(\$1626_t\); default_zero(\$v3743\); 
          default_zero(\$v3843\); default_zero(\$1220\); 
          default_zero(\$1638_x\); default_zero(\$v3746\); 
          default_zero(\$1298_i\); default_zero(\$v3627\); 
          default_zero(\$v2989\); default_zero(\$1327\); 
          default_zero(\$1203\); default_zero(\$911_i\); 
          default_zero(\$v3541\); default_zero(\$1307_i\); 
          default_zero(\$v3527\); default_zero(\$1315\); 
          default_zero(\$1426_t\); default_zero(\$v3450\); 
          default_zero(\$v3472\); default_zero(\$1678\); 
          default_zero(\$v3898\); default_zero(\$v3688\); 
          default_zero(\$v3643\); default_zero(\$v3607\); 
          default_zero(\$v3667\); default_zero(\$v3883\); 
          default_zero(\$1294\); default_zero(\$1500\); 
          default_zero(\$1603\); default_zero(\$v3874\); 
          default_zero(\$1423_print_value6133369_arg\); 
          default_zero(\$v3953\); default_zero(\$1164\); 
          default_zero(\$v3640\); default_zero(\$v3523\); 
          default_zero(\$1623\); default_zero(\$v3978\); 
          default_zero(\$v3752\); default_zero(\$1529\); 
          default_zero(\$1250\); default_zero(\$v3705\); 
          default_zero(\$v3702\); default_zero(\$1503\); 
          default_zero(\$1521_i\); default_zero(\$v3605\); 
          default_zero(\$1336\); default_zero(\$v3963\); 
          default_zero(\$1194\); default_zero(\$v3659\); 
          default_zero(\$v3714\); default_zero(\$v3500\); 
          default_zero(\$v3598\); default_zero(\$1446_t\); 
          default_zero(\$v3412\); default_zero(\$1625\); 
          default_zero(\$1073_loop667_arg\); default_zero(\$1285\); 
          default_zero(\$v3754\); default_zero(\$1504_i\); 
          default_zero(\$v3434\); default_zero(\$v3824\); 
          default_zero(\$1464_loop6693373_arg\); default_zero(\$v4025\); 
          default_zero(\$v3944\); default_zero(\$v3866\); 
          default_zero(\$1186_i\); default_zero(\$v3781\); 
          default_zero(\$v3464\); default_zero(\$v3709\); 
          default_zero(\$1519\); default_zero(\$v3804\); 
          default_zero(\$1541\); default_zero(\$v3873\); 
          default_zero(\$1464_loop6693373_result\); default_zero(\$v3700\); 
          default_zero(\$v2972\); default_zero(\$v4009\); 
          default_zero(\$v2916\); default_zero(\$v3949\); 
          default_zero(\$v3730\); default_zero(\$v1694\); 
          default_zero(\$v1666\); default_zero(\$1204_t\); 
          default_zero(\$411_show_rib6323359_result\); default_zero(\$1383\); 
          default_zero(\$v3690\); default_zero(\$v3830\); 
          default_zero(\$1158\); default_zero(\$1325\); 
          default_zero(\$v3780\); default_zero(\$v3482\); 
          default_zero(\$v3442\); default_zero(\$v3712\); 
          default_zero(\$1242_i\); default_zero(\$v3745\); 
          default_zero(\$v3787\); default_zero(\$v3853\); 
          default_zero(\$v3645\); default_zero(\$1053_i\); 
          default_zero(\$1108\); default_zero(\$v3985\); 
          default_zero(\$1584\); default_zero(\$v3943\); 
          default_zero(\$v3459\); default_zero(\$1109_i\); 
          default_zero(\$v3496\); default_zero(\$1577\); 
          default_zero(\$v3486\); default_zero(\$1680_i\); 
          default_zero(\$1009_t\); default_zero(\$v3839\); 
          default_zero(\$v3799\); default_zero(\$v3835\); 
          default_zero(\$v3771\); default_zero(\$v3964\); 
          default_zero(\$1511\); default_zero(\$v3542\); 
          default_zero(\$v3418\); default_zero(\$v3419\); 
          default_zero(\$411_show_rib6323357_result\); 
          default_zero(\$v3608\); default_zero(\$v3747\); 
          default_zero(\$v3719\); default_zero(\$v3692\); 
          default_zero(\$v3597\); default_zero(\$v3911\); 
          default_zero(\$v3591\); default_zero(\$v3869\); 
          default_zero(\$1277_i\); default_zero(\$v3860\); 
          default_zero(\$v3594\); default_zero(\$1651\); 
          default_zero(\$v3650\); default_zero(\$v3673\); 
          default_zero(\$1382\); default_zero(result3406); 
          default_zero(\$v3725\); default_zero(\$v3984\); 
          default_zero(\$v3798\); default_zero(\$1101_car\); 
          default_zero(\$v3704\); default_zero(\$v3681\); 
          default_zero(\$v3564\); default_zero(\$v3644\); 
          default_zero(\$v3919\); default_zero(\$1127\); 
          default_zero(\$v3759\); default_zero(\$1443\); 
          default_zero(\$v3983\); default_zero(\$1102\); 
          default_zero(\$1571_i\); default_zero(\$1259\); 
          default_zero(\$v4033\); default_zero(\$v3430\); 
          default_zero(\$v4001\); default_zero(\$v3578\); 
          default_zero(\$v3854\); default_zero(\$1107\); 
          default_zero(\$1673\); default_zero(\$1539\); 
          default_zero(\$v3711\); default_zero(\$v3593\); 
          default_zero(\$v3668\); default_zero(\$v2925\); 
          default_zero(\$1117\); default_zero(\$v3885\); 
          default_zero(\$1070_get_int640_arg\); default_zero(\$1183\); 
          default_zero(\$v2985\); default_zero(\$v3492\); 
          default_zero(\$1165_i\); default_zero(\$1656\); 
          default_zero(\$v3628\); default_zero(\$1384_i\); 
          default_zero(\$v4029\); default_zero(\$v3976\); 
          default_zero(\$1260_t\); default_zero(\$v3675\); 
          default_zero(\$v3961\); default_zero(\$1139_i\); 
          default_zero(\$v3731\); default_zero(\$1147\); 
          default_zero(\$1445\); default_zero(\$v3691\); 
          default_zero(\$v3931\); default_zero(\$v3858\); 
          default_zero(\$v3918\); default_zero(\$1049_i\); 
          default_zero(\$v3618\); default_zero(\$v2929\); 
          default_zero(\$v3467\); default_zero(\$1422\); 
          default_zero(\$v3875\); default_zero(\$v3825\); 
          default_zero(\$v3554\); default_zero(\$v3533\); 
          default_zero(\$1658\); default_zero(\$1653_c\); 
          default_zero(\$v3515\); default_zero(\$1492\); 
          default_zero(\$v3822\); default_zero(\$v3935\); 
          default_zero(\$v3726\); default_zero(\$v3755\); 
          default_zero(\$1655\); default_zero(\$v3716\); 
          default_zero(\$v4005\); default_zero(\$v3577\); 
          default_zero(\$1454_t\); default_zero(\$v3680\); 
          default_zero(\$v3572\); default_zero(\$1269_car\); 
          default_zero(\$1604\); default_zero(\$v3596\); 
          default_zero(\$v3905\); default_zero(\$1485\); 
          default_zero(\$v3570\); default_zero(\$v3620\); 
          default_zero(\$v3655\); default_zero(rdy3407); 
          default_zero(\$v3997\); default_zero(\$v3583\); 
          default_zero(\$v2976\); default_zero(\$1156\); 
          default_zero(\$1130_i\); default_zero(\$v3411\); 
          default_zero(\$v3488\); default_zero(\$v3831\); 
          default_zero(\$v3777\); default_zero(\$v3699\); 
          default_zero(\$v4021\); default_zero(\$v3689\); 
          default_zero(\$v3701\); default_zero(\$v3478\); 
          default_zero(\$1316_t\); default_zero(\$914\); 
          default_zero(\$v1704\); default_zero(\$v3848\); 
          default_zero(\$v3573\); default_zero(\$v3619\); 
          default_zero(\$v3887\); default_zero(\$v3765\); 
          default_zero(\$v3840\); default_zero(\$1490\); 
          default_zero(\$v3663\); default_zero(\$1444\); 
          default_zero(\$v3672\); default_zero(\$1605_i\); 
          default_zero(\$v3897\); default_zero(\$1270\); 
          default_zero(\$1230_t\); default_zero(\$1477_t\); 
          default_zero(\$1414_t\); default_zero(\$v3710\); 
          default_zero(\$1550\); default_zero(\$v3766\); 
          default_zero(\$1677\); default_zero(\$v3884\); 
          default_zero(\$v3579\); default_zero(\$v3409\); 
          default_zero(\$v3910\); default_zero(\$1491\); 
          default_zero(\$v3425\); default_zero(\$v3879\); 
          default_zero(\$v3465\); default_zero(\$v3625\); 
          default_zero(\$v3970\); default_zero(\$1157_car\); 
          default_zero(\$v3728\); default_zero(\$v3975\); 
          default_zero(\$v3556\); default_zero(\$v3410\); 
          default_zero(\$1396_i\); default_zero(\$v3847\); 
          default_zero(\$v3751\); default_zero(\$v3957\); 
          default_zero(\$1585\); default_zero(\$v3557\); 
          default_zero(\$1657\); default_zero(\$v3917\); 
          default_zero(\$v3633\); default_zero(\$v1713\); 
          default_zero(\$v3772\); default_zero(\$913\); 
          default_zero(\$1072_rest_loop668_arg\); default_zero(\$1428_i\); 
          default_zero(\$v3791\); default_zero(\$v3892\); 
          default_zero(\$1622\); default_zero(\$v3528\); 
          default_zero(\$v3481\); default_zero(\$v3909\); 
          default_zero(\$v3634\); default_zero(\$v3968\); 
          default_zero(\$1588_i\); default_zero(\$v3604\); 
          default_zero(\$v3829\); default_zero(\$v3760\); 
          default_zero(\$v3558\); default_zero(\$v3503\); 
          default_zero(\$v3501\); default_zero(\$1538\); 
          default_zero(\$v3841\); default_zero(\$1530_t\); 
          default_zero(\$v3649\); default_zero(\$v3563\); 
          default_zero(\$v3977\); default_zero(\$v3537\); 
          default_zero(\$1328\); default_zero(\$1587\); 
          default_zero(\$v3939\); default_zero(\$v3817\); 
          default_zero(\$v3809\); default_zero(\$411_show_rib6323359_arg\); 
          default_zero(\$v3727\); default_zero(\$1494\); 
          default_zero(\$1333\); default_zero(\$1393\); 
          default_zero(\$1214\); default_zero(\$v3785\); 
          default_zero(\$v3859\); default_zero(\$1138\); 
          default_zero(\$v3546\); default_zero(\$1276\); 
          default_zero(\$1163\); default_zero(\$v2950\); 
          default_zero(\$v3511\); default_zero(\$v3302\); 
          default_zero(\$v3732\); default_zero(\$v3982\); 
          default_zero(\$1595\); default_zero(\$v3865\); 
          default_zero(\$v3805\); default_zero(\$v1723\); 
          default_zero(\$v2920\); default_zero(\$v3315\); 
          default_zero(\$v3519\); default_zero(\$1306\); 
          default_zero(\$v3720\); default_zero(\$v402\); 
          default_zero(\$v3713\); default_zero(\$v3595\); 
          default_zero(\$1439\); default_zero(\$1438_k\); 
          default_zero(\$v3796\); default_zero(\$v3737\); 
          default_zero(\$1251_i\); default_zero(\$v3592\); 
          default_zero(\$v3868\); default_zero(\$v3971\); 
          default_zero(\$v3466\); default_zero(\$v3724\); 
          default_zero(\$v3761\); default_zero(\$1429_t\); 
          default_zero(\$v3642\); default_zero(\$v3473\); 
          default_zero(\$v3626\); default_zero(\$1542_t\); 
          default_zero(\$v3617\); default_zero(\$1395\); 
          default_zero(\$v3902\); default_zero(\$v3904\); 
          default_zero(\$v3742\); default_zero(\$v3550\); 
          default_zero(\$v3810\); default_zero(\$v3770\); 
          default_zero(\$1371_show_rib6323365_arg\); default_zero(\$1650\); 
          default_zero(\$v3816\); default_zero(\$v1675\); 
          default_zero(\$1520\); default_zero(\$1463\); 
          default_zero(\$1118_t\); default_zero(\$1467_tag\); 
          default_zero(\$v3803\); default_zero(\$1486\); 
          default_zero(\$v3568\); default_zero(\$v3471\); 
          default_zero(\$v3729\); default_zero(\$v3695\); 
          default_zero(\$v3989\); 
          default_zero(\$1371_show_rib6323365_result\); 
          default_zero(\$v3477\); default_zero(\$v3821\); 
          default_zero(\$v3786\); default_zero(\$v3636\); 
          default_zero(\$v3797\); default_zero(\$1148_t\); 
          default_zero(\$1239\); default_zero(\$1688\); 
          default_zero(\$v3927\); default_zero(\$v3815\); 
          default_zero(\$1126\); default_zero(\$v3823\); 
          default_zero(\$1182\); default_zero(\$v3641\); 
          default_zero(\$v3674\); default_zero(\$1501\); 
          default_zero(\$1213_car\); 
          default_zero(\$1423_print_value6133369_result\); 
          default_zero(\$v3849\); default_zero(\$1212\); 
          default_zero(\$1394\); default_zero(\$v3717\); 
          default_zero(\$v3679\); default_zero(\$1551\); 
          default_zero(\$v3694\); default_zero(\$v3606\); 
          default_zero(\$v3923\); default_zero(\$1569\); 
          default_zero(\$v3599\); default_zero(\$v3693\); 
          default_zero(\$1648_x\); default_zero(\$v3463\); 
          default_zero(\$v3738\); default_zero(\$v3502\); 
          default_zero(\$1275\); default_zero(\$v3416\); 
          default_zero(\$1614_t\); default_zero(\$v3903\); 
          default_zero(\$v3479\); default_zero(\$v3744\); 
          default_zero(\$1229\); default_zero(\$v3651\); 
          default_zero(\$v3814\); default_zero(\$1575\); 
          default_zero(\$v3945\); default_zero(\$1238\); 
          default_zero(\$1665\); default_zero(\$v4013\); 
          default_zero(\$v3893\); default_zero(\$v3867\); 
          default_zero(\$v3687\); default_zero(\$v3609\); 
          default_zero(\$v3736\); default_zero(\$v3635\); 
          default_zero(\$v3424\); default_zero(\$1404\); 
          default_zero(\$1570\); default_zero(\$v3417\); 
          default_zero(\$v3715\); default_zero(\$v3532\); 
          default_zero(\$v3886\); default_zero(\$v3773\); 
          default_zero(\$v3426\); default_zero(\$v3507\); 
          default_zero(\$v3778\); default_zero(\$v3569\); 
          default_zero(\$v3420\); default_zero(\$v3962\); 
          default_zero(\$v1685\); default_zero(\$1634\); 
          default_zero(\$1690\); default_zero(\$1295\); 
          default_zero(\$411_show_rib6323357_arg\); default_zero(\$v3480\); 
          default_zero(\$v4017\); 
          rdy <= "1";
          rdy3407 := "0";
          \state\ <= compute3408;
          
        else if run = '1' then
          case \state\ is
          when \$1069_list_tail637\ =>
            \$v3425\ := eclat_eq("00000000000000000000000000000000" & \$1069_list_tail637_arg\(32 to 63));
            if \$v3425\(0) = '1' then
              \$v3409\ := \$1069_list_tail637_arg\(0 to 31);
              
              \state\ <= \$1069_list_tail637\;
            else
              \$v3424\ := \$arr3399_ptr_take\;
              if \$v3424\(0) = '1' then
                \state\ <= q_wait3423;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1069_list_tail637_arg\(0 to 31)));
                \state\ <= pause_getI3421;
              end if;
            end if;
          when \$1070_get_int640\ =>
            \$v3442\ := \$arr3403_ptr_take\;
            if \$v3442\(0) = '1' then
              \state\ <= q_wait3441;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr\ <= 0;
              \state\ <= pause_getI3439;
            end if;
          when \$1072_rest_loop668\ =>
            \$v3533\ := eclat_lt("00000000000000000000000000000000" & \$1072_rest_loop668_arg\(36 to 67));
            if \$v3533\(0) = '1' then
              \$v3500\ := \$arr3400_ptr_take\;
              if \$v3500\(0) = '1' then
                \state\ <= q_wait3499;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr\ <= 0;
                \state\ <= pause_getI3497;
              end if;
            else
              \$v3532\ := \$arr3400_ptr_take\;
              if \$v3532\(0) = '1' then
                \state\ <= q_wait3531;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr\ <= 0;
                \state\ <= pause_getI3529;
              end if;
            end if;
          when \$1073_loop667\ =>
            \$v3747\ := eclat_lt("00000000000000000000000000000000" & \$1073_loop667_arg\(0 to 31));
            if \$v3747\(0) = '1' then
              \$v3591\ := \$arr3400_ptr_take\;
              if \$v3591\(0) = '1' then
                \state\ <= q_wait3590;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr\ <= 0;
                \state\ <= pause_getI3588;
              end if;
            else
              \$v3745\ := \$1073_loop667_arg\(68 to 103);
              \$v3746\ := \$v3745\(0 to 3);
              \$v3744\ := \$v3745\(4 to 35);
              case \$v3746\ is
              when "0010" =>
                \$1437\ := eclat_true;
                \$v3743\ := \$1437\;
                if \$v3743\(0) = '1' then
                  \$v3663\ := \$arr3399_ptr_take\;
                  if \$v3663\(0) = '1' then
                    \state\ <= q_wait3662;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                    \state\ <= pause_getI3660;
                  end if;
                else
                  \$v3742\ := \$arr3400_ptr_take\;
                  if \$v3742\(0) = '1' then
                    \state\ <= q_wait3741;
                  else
                    \$arr3400_ptr_take\(0) := '1';
                    \$arr3400_ptr\ <= 0;
                    \state\ <= pause_getI3739;
                  end if;
                end if;
              when others =>
                \$1437\ := eclat_false;
                \$v3743\ := \$1437\;
                if \$v3743\(0) = '1' then
                  \$v3663\ := \$arr3399_ptr_take\;
                  if \$v3663\(0) = '1' then
                    \state\ <= q_wait3662;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                    \state\ <= pause_getI3660;
                  end if;
                else
                  \$v3742\ := \$arr3400_ptr_take\;
                  if \$v3742\(0) = '1' then
                    \state\ <= q_wait3741;
                  else
                    \$arr3400_ptr_take\(0) := '1';
                    \$arr3400_ptr\ <= 0;
                    \state\ <= pause_getI3739;
                  end if;
                end if;
              end case;
            end if;
          when \$1113_forever6893378\ =>
            \state\ <= \$1113_forever6893378\;
          when \$1122_forever6893379\ =>
            \state\ <= \$1122_forever6893379\;
          when \$1134_forever6893380\ =>
            \state\ <= \$1134_forever6893380\;
          when \$1143_forever6893381\ =>
            \state\ <= \$1143_forever6893381\;
          when \$1152_forever6893382\ =>
            \state\ <= \$1152_forever6893382\;
          when \$1169_forever6893383\ =>
            \state\ <= \$1169_forever6893383\;
          when \$1178_forever6893384\ =>
            \state\ <= \$1178_forever6893384\;
          when \$1190_forever6893385\ =>
            \state\ <= \$1190_forever6893385\;
          when \$1199_forever6893386\ =>
            \state\ <= \$1199_forever6893386\;
          when \$1208_forever6893387\ =>
            \state\ <= \$1208_forever6893387\;
          when \$1225_forever6893388\ =>
            \state\ <= \$1225_forever6893388\;
          when \$1234_forever6893389\ =>
            \state\ <= \$1234_forever6893389\;
          when \$1246_forever6893390\ =>
            \state\ <= \$1246_forever6893390\;
          when \$1255_forever6893391\ =>
            \state\ <= \$1255_forever6893391\;
          when \$1264_forever6893392\ =>
            \state\ <= \$1264_forever6893392\;
          when \$1281_forever6893393\ =>
            \state\ <= \$1281_forever6893393\;
          when \$1290_forever6893394\ =>
            \state\ <= \$1290_forever6893394\;
          when \$1302_forever6893395\ =>
            \state\ <= \$1302_forever6893395\;
          when \$1311_forever6893396\ =>
            \state\ <= \$1311_forever6893396\;
          when \$1320_forever6893397\ =>
            \state\ <= \$1320_forever6893397\;
          when \$1371_show_rib6323365\ =>
            \$v3609\ := eclat_gt(\$1371_show_rib6323365_arg\(68 to 99) & \$1371_show_rib6323365_arg\(36 to 67));
            if \$v3609\(0) = '1' then
              \$v3597\ := \$1371_show_rib6323365_arg\(0 to 35);
              \$v3598\ := \$v3597\(0 to 3);
              \$v3596\ := \$v3597\(4 to 35);
              case \$v3598\ is
              when "0010" =>
                \$1382\ := eclat_true;
                \$v3595\ := \$1382\;
                if \$v3595\(0) = '1' then
                  \$1371_show_rib6323365_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \state\ <= \$1073_loop667\;
                else
                  \$v3593\ := \$1371_show_rib6323365_arg\(0 to 35);
                  \$v3594\ := \$v3593\(0 to 3);
                  \$v3592\ := \$v3593\(4 to 35);
                  case \$v3594\ is
                  when "0001" =>
                    \$1384_i\ := \$v3592\(0 to 31);
                    \$1383\ := \$1384_i\;
                    \$1371_show_rib6323365_result\ := eclat_unit;
                    eclat_print_int(\$1383\);
                    
                    \state\ <= \$1073_loop667\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$1388_forever6893337\;
                  end case;
                end if;
              when others =>
                \$1382\ := eclat_false;
                \$v3595\ := \$1382\;
                if \$v3595\(0) = '1' then
                  \$1371_show_rib6323365_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \state\ <= \$1073_loop667\;
                else
                  \$v3593\ := \$1371_show_rib6323365_arg\(0 to 35);
                  \$v3594\ := \$v3593\(0 to 3);
                  \$v3592\ := \$v3593\(4 to 35);
                  case \$v3594\ is
                  when "0001" =>
                    \$1384_i\ := \$v3592\(0 to 31);
                    \$1383\ := \$1384_i\;
                    \$1371_show_rib6323365_result\ := eclat_unit;
                    eclat_print_int(\$1383\);
                    
                    \state\ <= \$1073_loop667\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$1388_forever6893337\;
                  end case;
                end if;
              end case;
            else
              \$v3607\ := \$1371_show_rib6323365_arg\(0 to 35);
              \$v3608\ := \$v3607\(0 to 3);
              \$v3599\ := \$v3607\(4 to 35);
              case \$v3608\ is
              when "0000" =>
                \$1371_show_rib6323365_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \state\ <= \$1073_loop667\;
              when "0001" =>
                \$1380_i\ := \$v3599\(0 to 31);
                \$1371_show_rib6323365_result\ := eclat_unit;
                eclat_print_int(\$1380_i\);
                
                \state\ <= \$1073_loop667\;
              when "0010" =>
                \$v3605\ := \$1371_show_rib6323365_arg\(0 to 35);
                \$v3606\ := \$v3605\(0 to 3);
                \$v3600\ := \$v3605\(4 to 35);
                case \$v3606\ is
                when "0010" =>
                  \$1049_i\ := \$v3600\(0 to 31);
                  \$v3604\ := \$arr3399_ptr_take\;
                  if \$v3604\(0) = '1' then
                    \state\ <= q_wait3603;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
                    \state\ <= pause_getI3601;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$373_forever6893336\;
                end case;
              when others =>
                
              end case;
            end if;
          when \$1388_forever6893337\ =>
            \state\ <= \$1388_forever6893337\;
          when \$1400_forever6893366\ =>
            \state\ <= \$1400_forever6893366\;
          when \$1410_forever6893367\ =>
            \state\ <= \$1410_forever6893367\;
          when \$1418_forever6893368\ =>
            \state\ <= \$1418_forever6893368\;
          when \$1423_print_value6133369\ =>
            \$v3643\ := \$1423_print_value6133369_arg\;
            \$v3644\ := \$v3643\(0 to 3);
            \$v3635\ := \$v3643\(4 to 35);
            case \$v3644\ is
            when "0010" =>
              \$1426_t\ := \$v3635\(0 to 31);
              \$v3641\ := "0010" & \$1426_t\;
              \$v3642\ := \$v3641\(0 to 3);
              \$v3636\ := \$v3641\(4 to 35);
              case \$v3642\ is
              when "0010" =>
                \$1049_i\ := \$v3636\(0 to 31);
                \$v3640\ := \$arr3399_ptr_take\;
                if \$v3640\(0) = '1' then
                  \state\ <= q_wait3639;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
                  \state\ <= pause_getI3637;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_rib expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$373_forever6893335\;
              end case;
            when "0000" =>
              \$1423_print_value6133369_result\ := eclat_unit;
              eclat_print_string(of_string("Nil"));
              
              eclat_print_string(of_string("printed tag dfe code\n"));
              
              \$v3633\ := \$1073_loop667_arg\(104 to 139);
              \$v3634\ := \$v3633\(0 to 3);
              \$v3628\ := \$v3633\(4 to 35);
              case \$v3634\ is
              when "0010" =>
                \$1414_t\ := \$v3628\(0 to 31);
                \$v3632\ := \$arr3399_ptr_take\;
                if \$v3632\(0) = '1' then
                  \state\ <= q_wait3631;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1414_t\));
                  \state\ <= pause_getI3629;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_tag_triplet expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1418_forever6893368\;
              end case;
            when "0001" =>
              \$1428_i\ := \$v3635\(0 to 31);
              \$1423_print_value6133369_result\ := eclat_unit;
              eclat_print_int(\$1428_i\);
              
              eclat_print_string(of_string("printed tag dfe code\n"));
              
              \$v3633\ := \$1073_loop667_arg\(104 to 139);
              \$v3634\ := \$v3633\(0 to 3);
              \$v3628\ := \$v3633\(4 to 35);
              case \$v3634\ is
              when "0010" =>
                \$1414_t\ := \$v3628\(0 to 31);
                \$v3632\ := \$arr3399_ptr_take\;
                if \$v3632\(0) = '1' then
                  \state\ <= q_wait3631;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1414_t\));
                  \state\ <= pause_getI3629;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_tag_triplet expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1418_forever6893368\;
              end case;
            when others =>
              
            end case;
          when \$1433_forever6893370\ =>
            \state\ <= \$1433_forever6893370\;
          when \$1450_forever6893371\ =>
            \state\ <= \$1450_forever6893371\;
          when \$1458_forever6893372\ =>
            \state\ <= \$1458_forever6893372\;
          when \$1464_loop6693373\ =>
            \$v3737\ := \$1464_loop6693373_arg\;
            \$v3738\ := \$v3737\(0 to 3);
            \$v3732\ := \$v3737\(4 to 35);
            case \$v3738\ is
            when "0010" =>
              \$1477_t\ := \$v3732\(0 to 31);
              \$v3736\ := \$arr3399_ptr_take\;
              if \$v3736\(0) = '1' then
                \state\ <= q_wait3735;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1477_t\));
                \state\ <= pause_getI3733;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1481_forever6893360\;
            end case;
          when \$1473_forever6893356\ =>
            \state\ <= \$1473_forever6893356\;
          when \$1481_forever6893360\ =>
            \state\ <= \$1481_forever6893360\;
          when \$1515_forever6893374\ =>
            \state\ <= \$1515_forever6893374\;
          when \$1525_forever6893375\ =>
            \state\ <= \$1525_forever6893375\;
          when \$1534_forever6893376\ =>
            \state\ <= \$1534_forever6893376\;
          when \$1546_forever6893377\ =>
            \state\ <= \$1546_forever6893377\;
          when \$1599_forever6893361\ =>
            \state\ <= \$1599_forever6893361\;
          when \$1609_forever6893362\ =>
            \state\ <= \$1609_forever6893362\;
          when \$1618_forever6893363\ =>
            \state\ <= \$1618_forever6893363\;
          when \$1630_forever6893364\ =>
            \state\ <= \$1630_forever6893364\;
          when \$1669_forever6893338\ =>
            \state\ <= \$1669_forever6893338\;
          when \$1684_forever6893339\ =>
            \state\ <= \$1684_forever6893339\;
          when \$373_forever6893335\ =>
            \state\ <= \$373_forever6893335\;
          when \$373_forever6893336\ =>
            \state\ <= \$373_forever6893336\;
          when \$373_forever6893337\ =>
            \state\ <= \$373_forever6893337\;
          when \$373_forever6893358\ =>
            \state\ <= \$373_forever6893358\;
          when \$411_show_rib6323357\ =>
            \$v3704\ := eclat_gt(\$411_show_rib6323357_arg\(68 to 99) & \$411_show_rib6323357_arg\(36 to 67));
            if \$v3704\(0) = '1' then
              \$v3692\ := \$411_show_rib6323357_arg\(0 to 35);
              \$v3693\ := \$v3692\(0 to 3);
              \$v3691\ := \$v3692\(4 to 35);
              case \$v3693\ is
              when "0010" =>
                \$913\ := eclat_true;
                \$v3690\ := \$913\;
                if \$v3690\(0) = '1' then
                  \$411_show_rib6323357_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                  \$1438_k\ := \$1464_loop6693373_result\;
                  \$v3685\ := \$arr3399_ptr_take\;
                  if \$v3685\(0) = '1' then
                    \state\ <= q_wait3684;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                    \state\ <= pause_getI3682;
                  end if;
                else
                  \$v3688\ := \$411_show_rib6323357_arg\(0 to 35);
                  \$v3689\ := \$v3688\(0 to 3);
                  \$v3687\ := \$v3688\(4 to 35);
                  case \$v3689\ is
                  when "0001" =>
                    \$1053_i\ := \$v3687\(0 to 31);
                    \$914\ := \$1053_i\;
                    \$411_show_rib6323357_result\ := eclat_unit;
                    eclat_print_int(\$914\);
                    
                    \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                    \$1438_k\ := \$1464_loop6693373_result\;
                    \$v3685\ := \$arr3399_ptr_take\;
                    if \$v3685\(0) = '1' then
                      \state\ <= q_wait3684;
                    else
                      \$arr3399_ptr_take\(0) := '1';
                      \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                      \state\ <= pause_getI3682;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893337\;
                  end case;
                end if;
              when others =>
                \$913\ := eclat_false;
                \$v3690\ := \$913\;
                if \$v3690\(0) = '1' then
                  \$411_show_rib6323357_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                  \$1438_k\ := \$1464_loop6693373_result\;
                  \$v3685\ := \$arr3399_ptr_take\;
                  if \$v3685\(0) = '1' then
                    \state\ <= q_wait3684;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                    \state\ <= pause_getI3682;
                  end if;
                else
                  \$v3688\ := \$411_show_rib6323357_arg\(0 to 35);
                  \$v3689\ := \$v3688\(0 to 3);
                  \$v3687\ := \$v3688\(4 to 35);
                  case \$v3689\ is
                  when "0001" =>
                    \$1053_i\ := \$v3687\(0 to 31);
                    \$914\ := \$1053_i\;
                    \$411_show_rib6323357_result\ := eclat_unit;
                    eclat_print_int(\$914\);
                    
                    \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                    \$1438_k\ := \$1464_loop6693373_result\;
                    \$v3685\ := \$arr3399_ptr_take\;
                    if \$v3685\(0) = '1' then
                      \state\ <= q_wait3684;
                    else
                      \$arr3399_ptr_take\(0) := '1';
                      \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                      \state\ <= pause_getI3682;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893337\;
                  end case;
                end if;
              end case;
            else
              \$v3702\ := \$411_show_rib6323357_arg\(0 to 35);
              \$v3703\ := \$v3702\(0 to 3);
              \$v3694\ := \$v3702\(4 to 35);
              case \$v3703\ is
              when "0000" =>
                \$411_show_rib6323357_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                \$1438_k\ := \$1464_loop6693373_result\;
                \$v3685\ := \$arr3399_ptr_take\;
                if \$v3685\(0) = '1' then
                  \state\ <= q_wait3684;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                  \state\ <= pause_getI3682;
                end if;
              when "0001" =>
                \$911_i\ := \$v3694\(0 to 31);
                \$411_show_rib6323357_result\ := eclat_unit;
                eclat_print_int(\$911_i\);
                
                \$1464_loop6693373_result\ := \$1464_loop6693373_arg\;
                \$1438_k\ := \$1464_loop6693373_result\;
                \$v3685\ := \$arr3399_ptr_take\;
                if \$v3685\(0) = '1' then
                  \state\ <= q_wait3684;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
                  \state\ <= pause_getI3682;
                end if;
              when "0010" =>
                \$v3700\ := \$411_show_rib6323357_arg\(0 to 35);
                \$v3701\ := \$v3700\(0 to 3);
                \$v3695\ := \$v3700\(4 to 35);
                case \$v3701\ is
                when "0010" =>
                  \$1049_i\ := \$v3695\(0 to 31);
                  \$v3699\ := \$arr3399_ptr_take\;
                  if \$v3699\(0) = '1' then
                    \state\ <= q_wait3698;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
                    \state\ <= pause_getI3696;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$373_forever6893336\;
                end case;
              when others =>
                
              end case;
            end if;
          when \$411_show_rib6323359\ =>
            \$v3729\ := eclat_gt(\$411_show_rib6323359_arg\(68 to 99) & \$411_show_rib6323359_arg\(36 to 67));
            if \$v3729\(0) = '1' then
              \$v3717\ := \$411_show_rib6323359_arg\(0 to 35);
              \$v3718\ := \$v3717\(0 to 3);
              \$v3716\ := \$v3717\(4 to 35);
              case \$v3718\ is
              when "0010" =>
                \$913\ := eclat_true;
                \$v3715\ := \$913\;
                if \$v3715\(0) = '1' then
                  \$411_show_rib6323359_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$v3710\ := \$1464_loop6693373_arg\;
                  \$v3711\ := \$v3710\(0 to 3);
                  \$v3705\ := \$v3710\(4 to 35);
                  case \$v3711\ is
                  when "0010" =>
                    \$1009_t\ := \$v3705\(0 to 31);
                    \$v3709\ := \$arr3399_ptr_take\;
                    if \$v3709\(0) = '1' then
                      \state\ <= q_wait3708;
                    else
                      \$arr3399_ptr_take\(0) := '1';
                      \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                      \state\ <= pause_getI3706;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893358\;
                  end case;
                else
                  \$v3713\ := \$411_show_rib6323359_arg\(0 to 35);
                  \$v3714\ := \$v3713\(0 to 3);
                  \$v3712\ := \$v3713\(4 to 35);
                  case \$v3714\ is
                  when "0001" =>
                    \$1053_i\ := \$v3712\(0 to 31);
                    \$914\ := \$1053_i\;
                    \$411_show_rib6323359_result\ := eclat_unit;
                    eclat_print_int(\$914\);
                    
                    \$v3710\ := \$1464_loop6693373_arg\;
                    \$v3711\ := \$v3710\(0 to 3);
                    \$v3705\ := \$v3710\(4 to 35);
                    case \$v3711\ is
                    when "0010" =>
                      \$1009_t\ := \$v3705\(0 to 31);
                      \$v3709\ := \$arr3399_ptr_take\;
                      if \$v3709\(0) = '1' then
                        \state\ <= q_wait3708;
                      else
                        \$arr3399_ptr_take\(0) := '1';
                        \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                        \state\ <= pause_getI3706;
                      end if;
                    when others =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \state\ <= \$373_forever6893358\;
                    end case;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893337\;
                  end case;
                end if;
              when others =>
                \$913\ := eclat_false;
                \$v3715\ := \$913\;
                if \$v3715\(0) = '1' then
                  \$411_show_rib6323359_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$v3710\ := \$1464_loop6693373_arg\;
                  \$v3711\ := \$v3710\(0 to 3);
                  \$v3705\ := \$v3710\(4 to 35);
                  case \$v3711\ is
                  when "0010" =>
                    \$1009_t\ := \$v3705\(0 to 31);
                    \$v3709\ := \$arr3399_ptr_take\;
                    if \$v3709\(0) = '1' then
                      \state\ <= q_wait3708;
                    else
                      \$arr3399_ptr_take\(0) := '1';
                      \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                      \state\ <= pause_getI3706;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893358\;
                  end case;
                else
                  \$v3713\ := \$411_show_rib6323359_arg\(0 to 35);
                  \$v3714\ := \$v3713\(0 to 3);
                  \$v3712\ := \$v3713\(4 to 35);
                  case \$v3714\ is
                  when "0001" =>
                    \$1053_i\ := \$v3712\(0 to 31);
                    \$914\ := \$1053_i\;
                    \$411_show_rib6323359_result\ := eclat_unit;
                    eclat_print_int(\$914\);
                    
                    \$v3710\ := \$1464_loop6693373_arg\;
                    \$v3711\ := \$v3710\(0 to 3);
                    \$v3705\ := \$v3710\(4 to 35);
                    case \$v3711\ is
                    when "0010" =>
                      \$1009_t\ := \$v3705\(0 to 31);
                      \$v3709\ := \$arr3399_ptr_take\;
                      if \$v3709\(0) = '1' then
                        \state\ <= q_wait3708;
                      else
                        \$arr3399_ptr_take\(0) := '1';
                        \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                        \state\ <= pause_getI3706;
                      end if;
                    when others =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \state\ <= \$373_forever6893358\;
                    end case;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$373_forever6893337\;
                  end case;
                end if;
              end case;
            else
              \$v3727\ := \$411_show_rib6323359_arg\(0 to 35);
              \$v3728\ := \$v3727\(0 to 3);
              \$v3719\ := \$v3727\(4 to 35);
              case \$v3728\ is
              when "0000" =>
                \$411_show_rib6323359_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \$v3710\ := \$1464_loop6693373_arg\;
                \$v3711\ := \$v3710\(0 to 3);
                \$v3705\ := \$v3710\(4 to 35);
                case \$v3711\ is
                when "0010" =>
                  \$1009_t\ := \$v3705\(0 to 31);
                  \$v3709\ := \$arr3399_ptr_take\;
                  if \$v3709\(0) = '1' then
                    \state\ <= q_wait3708;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                    \state\ <= pause_getI3706;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$373_forever6893358\;
                end case;
              when "0001" =>
                \$911_i\ := \$v3719\(0 to 31);
                \$411_show_rib6323359_result\ := eclat_unit;
                eclat_print_int(\$911_i\);
                
                \$v3710\ := \$1464_loop6693373_arg\;
                \$v3711\ := \$v3710\(0 to 3);
                \$v3705\ := \$v3710\(4 to 35);
                case \$v3711\ is
                when "0010" =>
                  \$1009_t\ := \$v3705\(0 to 31);
                  \$v3709\ := \$arr3399_ptr_take\;
                  if \$v3709\(0) = '1' then
                    \state\ <= q_wait3708;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
                    \state\ <= pause_getI3706;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$373_forever6893358\;
                end case;
              when "0010" =>
                \$v3725\ := \$411_show_rib6323359_arg\(0 to 35);
                \$v3726\ := \$v3725\(0 to 3);
                \$v3720\ := \$v3725\(4 to 35);
                case \$v3726\ is
                when "0010" =>
                  \$1049_i\ := \$v3720\(0 to 31);
                  \$v3724\ := \$arr3399_ptr_take\;
                  if \$v3724\(0) = '1' then
                    \state\ <= q_wait3723;
                  else
                    \$arr3399_ptr_take\(0) := '1';
                    \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
                    \state\ <= pause_getI3721;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$373_forever6893336\;
                end case;
              when others =>
                
              end case;
            end if;
          when pause_getI3413 =>
            \state\ <= pause_getII3414;
          when pause_getI3421 =>
            \state\ <= pause_getII3422;
          when pause_getI3431 =>
            \state\ <= pause_getII3432;
          when pause_getI3435 =>
            \state\ <= pause_getII3436;
          when pause_getI3439 =>
            \state\ <= pause_getII3440;
          when pause_getI3443 =>
            \state\ <= pause_getII3444;
          when pause_getI3456 =>
            \state\ <= pause_getII3457;
          when pause_getI3468 =>
            \state\ <= pause_getII3469;
          when pause_getI3474 =>
            \state\ <= pause_getII3475;
          when pause_getI3483 =>
            \state\ <= pause_getII3484;
          when pause_getI3489 =>
            \state\ <= pause_getII3490;
          when pause_getI3493 =>
            \state\ <= pause_getII3494;
          when pause_getI3497 =>
            \state\ <= pause_getII3498;
          when pause_getI3512 =>
            \state\ <= pause_getII3513;
          when pause_getI3524 =>
            \state\ <= pause_getII3525;
          when pause_getI3529 =>
            \state\ <= pause_getII3530;
          when pause_getI3534 =>
            \state\ <= pause_getII3535;
          when pause_getI3547 =>
            \state\ <= pause_getII3548;
          when pause_getI3559 =>
            \state\ <= pause_getII3560;
          when pause_getI3565 =>
            \state\ <= pause_getII3566;
          when pause_getI3574 =>
            \state\ <= pause_getII3575;
          when pause_getI3580 =>
            \state\ <= pause_getII3581;
          when pause_getI3584 =>
            \state\ <= pause_getII3585;
          when pause_getI3588 =>
            \state\ <= pause_getII3589;
          when pause_getI3601 =>
            \state\ <= pause_getII3602;
          when pause_getI3610 =>
            \state\ <= pause_getII3611;
          when pause_getI3629 =>
            \state\ <= pause_getII3630;
          when pause_getI3637 =>
            \state\ <= pause_getII3638;
          when pause_getI3646 =>
            \state\ <= pause_getII3647;
          when pause_getI3656 =>
            \state\ <= pause_getII3657;
          when pause_getI3660 =>
            \state\ <= pause_getII3661;
          when pause_getI3669 =>
            \state\ <= pause_getII3670;
          when pause_getI3676 =>
            \state\ <= pause_getII3677;
          when pause_getI3682 =>
            \state\ <= pause_getII3683;
          when pause_getI3696 =>
            \state\ <= pause_getII3697;
          when pause_getI3706 =>
            \state\ <= pause_getII3707;
          when pause_getI3721 =>
            \state\ <= pause_getII3722;
          when pause_getI3733 =>
            \state\ <= pause_getII3734;
          when pause_getI3739 =>
            \state\ <= pause_getII3740;
          when pause_getI3756 =>
            \state\ <= pause_getII3757;
          when pause_getI3762 =>
            \state\ <= pause_getII3763;
          when pause_getI3774 =>
            \state\ <= pause_getII3775;
          when pause_getI3782 =>
            \state\ <= pause_getII3783;
          when pause_getI3788 =>
            \state\ <= pause_getII3789;
          when pause_getI3800 =>
            \state\ <= pause_getII3801;
          when pause_getI3806 =>
            \state\ <= pause_getII3807;
          when pause_getI3818 =>
            \state\ <= pause_getII3819;
          when pause_getI3826 =>
            \state\ <= pause_getII3827;
          when pause_getI3832 =>
            \state\ <= pause_getII3833;
          when pause_getI3844 =>
            \state\ <= pause_getII3845;
          when pause_getI3850 =>
            \state\ <= pause_getII3851;
          when pause_getI3862 =>
            \state\ <= pause_getII3863;
          when pause_getI3870 =>
            \state\ <= pause_getII3871;
          when pause_getI3876 =>
            \state\ <= pause_getII3877;
          when pause_getI3888 =>
            \state\ <= pause_getII3889;
          when pause_getI3894 =>
            \state\ <= pause_getII3895;
          when pause_getI3906 =>
            \state\ <= pause_getII3907;
          when pause_getI3914 =>
            \state\ <= pause_getII3915;
          when pause_getI3920 =>
            \state\ <= pause_getII3921;
          when pause_getI3928 =>
            \state\ <= pause_getII3929;
          when pause_getI3936 =>
            \state\ <= pause_getII3937;
          when pause_getI3946 =>
            \state\ <= pause_getII3947;
          when pause_getI3954 =>
            \state\ <= pause_getII3955;
          when pause_getII3414 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1673\ := \$arr3399_value\;
            \$v3411\ := \$1673\(36 to 71);
            \$v3412\ := \$v3411\(0 to 3);
            \$v3410\ := \$v3411\(4 to 35);
            case \$v3412\ is
            when "0010" =>
              \$1680_i\ := \$v3410\(0 to 31);
              \$1678\ := \$1680_i\;
              \$1677\ := \$1678\ & eclat_sub(\$1069_list_tail637_arg\(32 to 63) & "00000000000000000000000000000001");
              \$1069_list_tail637_arg\ := \$1677\;
              \state\ <= \$1069_list_tail637\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1684_forever6893339\;
            end case;
          when pause_getII3422 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1690\ := \$arr3399_value\;
            \$1688\ := \$1690\(36 to 71);
            \$v3419\ := \$1688\;
            \$v3420\ := \$v3419\(0 to 3);
            \$v3418\ := \$v3419\(4 to 35);
            case \$v3420\ is
            when "0010" =>
              \$1665\ := eclat_true;
              \$v3417\ := \$1665\;
              if \$v3417\(0) = '1' then
                \$v3416\ := \$arr3399_ptr_take\;
                if \$v3416\(0) = '1' then
                  \state\ <= q_wait3415;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1069_list_tail637_arg\(0 to 31)));
                  \state\ <= pause_getI3413;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("list_tail"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1669_forever6893338\;
              end if;
            when others =>
              \$1665\ := eclat_false;
              \$v3417\ := \$1665\;
              if \$v3417\(0) = '1' then
                \$v3416\ := \$arr3399_ptr_take\;
                if \$v3416\(0) = '1' then
                  \state\ <= q_wait3415;
                else
                  \$arr3399_ptr_take\(0) := '1';
                  \$arr3399_ptr\ <= to_integer(unsigned(\$1069_list_tail637_arg\(0 to 31)));
                  \state\ <= pause_getI3413;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("list_tail"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1669_forever6893338\;
              end if;
            end case;
          when pause_getII3432 =>
            \$arr3403_ptr_take\(0) := '0';
            \$1657\ := \$arr3403_value\;
            \$1656\ := \$1657\ & "00000000000000000000000000000001";
            \$1655\ := eclat_add(\$1656\);
            \$v3430\ := \$arr3403_ptr_take\;
            if \$v3430\(0) = '1' then
              \state\ <= q_wait3429;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr_write\ <= 0;
              \$arr3403_write_request\ <= '1';
              \$arr3403_write\ <= \$1655\;
              \state\ <= pause_setI3427;
            end if;
          when pause_getII3436 =>
            \$arr3398_ptr_take\(0) := '0';
            \$1653_c\ := \$arr3398_value\;
            \$v3434\ := \$arr3403_ptr_take\;
            if \$v3434\(0) = '1' then
              \state\ <= q_wait3433;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr\ <= 0;
              \state\ <= pause_getI3431;
            end if;
          when pause_getII3440 =>
            \$arr3403_ptr_take\(0) := '0';
            \$1658\ := \$arr3403_value\;
            \$v3438\ := \$arr3398_ptr_take\;
            if \$v3438\(0) = '1' then
              \state\ <= q_wait3437;
            else
              \$arr3398_ptr_take\(0) := '1';
              \$arr3398_ptr\ <= to_integer(unsigned(\$1658\));
              \state\ <= pause_getI3435;
            end if;
          when pause_getII3444 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1587\ := \$arr3404_value\;
            \$1585\ := "0010" & \$1587\;
            \$1584\ := \$1585\ & eclat_sub(\$1072_rest_loop668_arg\(36 to 67) & "00000000000000000000000000000001");
            \$1072_rest_loop668_arg\ := \$1584\ & \$1072_rest_loop668_arg\(68 to 99) & \$1072_rest_loop668_arg\(100 to 131);
            \state\ <= \$1072_rest_loop668\;
          when pause_getII3457 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1588_i\ := \$arr3404_value\;
            \$v3455\ := \$arr3399_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3451\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1588_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1578\(0 to 35) & \$1072_rest_loop668_arg\(0 to 35) & "0001" & \$v3451\;
              \state\ <= pause_setI3452;
            end if;
          when pause_getII3469 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2972\ := \$arr3399_value\;
            \$1604\ := \$v2972\(36 to 71);
            \$v3465\ := \$1604\;
            \$v3466\ := \$v3465\(0 to 3);
            \$v3464\ := \$v3465\(4 to 35);
            case \$v3466\ is
            when "0010" =>
              \$1605_i\ := \$v3464\(0 to 31);
              \$1603\ := \$1605_i\;
              \$v3463\ := \$arr3400_ptr_take\;
              if \$v3463\(0) = '1' then
                \state\ <= q_wait3462;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr_write\ <= 0;
                \$arr3400_write_request\ <= '1';
                \$arr3400_write\ <= \$1603\;
                \state\ <= pause_setI3460;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1609_forever6893362\;
            end case;
          when pause_getII3475 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1622\ := \$arr3400_value\;
            \$1613\ := "0010" & \$1622\;
            \$v3472\ := \$1613\;
            \$v3473\ := \$v3472\(0 to 3);
            \$v3467\ := \$v3472\(4 to 35);
            case \$v3473\ is
            when "0010" =>
              \$1614_t\ := \$v3467\(0 to 31);
              \$v3471\ := \$arr3399_ptr_take\;
              if \$v3471\(0) = '1' then
                \state\ <= q_wait3470;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1614_t\));
                \state\ <= pause_getI3468;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1618_forever6893363\;
            end case;
          when pause_getII3484 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2976\ := \$arr3399_value\;
            \$1623\ := \$v2976\(36 to 71);
            \$v3480\ := \$1623\;
            \$v3481\ := \$v3480\(0 to 3);
            \$v3479\ := \$v3480\(4 to 35);
            case \$v3481\ is
            when "0010" =>
              \$1595\ := eclat_true;
              \$v3478\ := \$1595\;
              if \$v3478\(0) = '1' then
                \$v3477\ := \$arr3400_ptr_take\;
                if \$v3477\(0) = '1' then
                  \state\ <= q_wait3476;
                else
                  \$arr3400_ptr_take\(0) := '1';
                  \$arr3400_ptr\ <= 0;
                  \state\ <= pause_getI3474;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1599_forever6893361\;
              end if;
            when others =>
              \$1595\ := eclat_false;
              \$v3478\ := \$1595\;
              if \$v3478\(0) = '1' then
                \$v3477\ := \$arr3400_ptr_take\;
                if \$v3477\(0) = '1' then
                  \state\ <= q_wait3476;
                else
                  \$arr3400_ptr_take\(0) := '1';
                  \$arr3400_ptr\ <= 0;
                  \state\ <= pause_getI3474;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1599_forever6893361\;
              end if;
            end case;
          when pause_getII3490 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1634\ := \$arr3400_value\;
            \$1625\ := "0010" & \$1634\;
            \$v3487\ := \$1625\;
            \$v3488\ := \$v3487\(0 to 3);
            \$v3482\ := \$v3487\(4 to 35);
            case \$v3488\ is
            when "0010" =>
              \$1626_t\ := \$v3482\(0 to 31);
              \$v3486\ := \$arr3399_ptr_take\;
              if \$v3486\(0) = '1' then
                \state\ <= q_wait3485;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1626_t\));
                \state\ <= pause_getI3483;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1630_forever6893364\;
            end case;
          when pause_getII3494 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1578\ := \$arr3399_value\;
            \$v3492\ := \$arr3400_ptr_take\;
            if \$v3492\(0) = '1' then
              \state\ <= q_wait3491;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3489;
            end if;
          when pause_getII3498 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1635\ := \$arr3400_value\;
            \$v3496\ := \$arr3399_ptr_take\;
            if \$v3496\(0) = '1' then
              \state\ <= q_wait3495;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1635\));
              \state\ <= pause_getI3493;
            end if;
          when pause_getII3513 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1569\ := \$arr3404_value\;
            \$v3511\ := \$arr3400_ptr_take\;
            if \$v3511\(0) = '1' then
              \state\ <= q_wait3510;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= \$1569\;
              \state\ <= pause_setI3508;
            end if;
          when pause_getII3525 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1571_i\ := \$arr3404_value\;
            \$v3523\ := \$arr3399_ptr_take\;
            if \$v3523\(0) = '1' then
              \state\ <= q_wait3522;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1571_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1570\;
              \state\ <= pause_setI3520;
            end if;
          when pause_getII3530 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1577\ := \$arr3400_value\;
            \$1575\ := "0010" & \$1577\;
            \$v3528\ := "00000000000000000000000000000000";
            \$1570\ := \$1072_rest_loop668_arg\(0 to 35) & \$1575\ & "0001" & \$v3528\;
            \$v3527\ := \$arr3404_ptr_take\;
            if \$v3527\(0) = '1' then
              \state\ <= q_wait3526;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3524;
            end if;
          when pause_getII3535 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1503\ := \$arr3404_value\;
            \$1501\ := "0010" & \$1503\;
            \$1500\ := eclat_sub(\$1073_loop667_arg\(0 to 31) & "00000000000000000000000000000001") & \$1501\;
            \$1073_loop667_arg\ := \$1500\ & \$1073_loop667_arg\(68 to 103) & \$1073_loop667_arg\(104 to 139) & \$1073_loop667_arg\(140 to 171);
            \state\ <= \$1073_loop667\;
          when pause_getII3548 =>
            \$arr3404_ptr_take\(0) := '0';
            \$1504_i\ := \$arr3404_value\;
            \$v3546\ := \$arr3399_ptr_take\;
            if \$v3546\(0) = '1' then
              \state\ <= q_wait3545;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3542\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1504_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1494\(0 to 35) & \$1073_loop667_arg\(32 to 67) & "0001" & \$v3542\;
              \state\ <= pause_setI3543;
            end if;
          when pause_getII3560 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2946\ := \$arr3399_value\;
            \$1520\ := \$v2946\(36 to 71);
            \$v3556\ := \$1520\;
            \$v3557\ := \$v3556\(0 to 3);
            \$v3555\ := \$v3556\(4 to 35);
            case \$v3557\ is
            when "0010" =>
              \$1521_i\ := \$v3555\(0 to 31);
              \$1519\ := \$1521_i\;
              \$v3554\ := \$arr3400_ptr_take\;
              if \$v3554\(0) = '1' then
                \state\ <= q_wait3553;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr_write\ <= 0;
                \$arr3400_write_request\ <= '1';
                \$arr3400_write\ <= \$1519\;
                \state\ <= pause_setI3551;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1525_forever6893375\;
            end case;
          when pause_getII3566 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1538\ := \$arr3400_value\;
            \$1529\ := "0010" & \$1538\;
            \$v3563\ := \$1529\;
            \$v3564\ := \$v3563\(0 to 3);
            \$v3558\ := \$v3563\(4 to 35);
            case \$v3564\ is
            when "0010" =>
              \$1530_t\ := \$v3558\(0 to 31);
              \$v3562\ := \$arr3399_ptr_take\;
              if \$v3562\(0) = '1' then
                \state\ <= q_wait3561;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1530_t\));
                \state\ <= pause_getI3559;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1534_forever6893376\;
            end case;
          when pause_getII3575 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2950\ := \$arr3399_value\;
            \$1539\ := \$v2950\(36 to 71);
            \$v3571\ := \$1539\;
            \$v3572\ := \$v3571\(0 to 3);
            \$v3570\ := \$v3571\(4 to 35);
            case \$v3572\ is
            when "0010" =>
              \$1511\ := eclat_true;
              \$v3569\ := \$1511\;
              if \$v3569\(0) = '1' then
                \$v3568\ := \$arr3400_ptr_take\;
                if \$v3568\(0) = '1' then
                  \state\ <= q_wait3567;
                else
                  \$arr3400_ptr_take\(0) := '1';
                  \$arr3400_ptr\ <= 0;
                  \state\ <= pause_getI3565;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1515_forever6893374\;
              end if;
            when others =>
              \$1511\ := eclat_false;
              \$v3569\ := \$1511\;
              if \$v3569\(0) = '1' then
                \$v3568\ := \$arr3400_ptr_take\;
                if \$v3568\(0) = '1' then
                  \state\ <= q_wait3567;
                else
                  \$arr3400_ptr_take\(0) := '1';
                  \$arr3400_ptr\ <= 0;
                  \state\ <= pause_getI3565;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1515_forever6893374\;
              end if;
            end case;
          when pause_getII3581 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1550\ := \$arr3400_value\;
            \$1541\ := "0010" & \$1550\;
            \$v3578\ := \$1541\;
            \$v3579\ := \$v3578\(0 to 3);
            \$v3573\ := \$v3578\(4 to 35);
            case \$v3579\ is
            when "0010" =>
              \$1542_t\ := \$v3573\(0 to 31);
              \$v3577\ := \$arr3399_ptr_take\;
              if \$v3577\(0) = '1' then
                \state\ <= q_wait3576;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1542_t\));
                \state\ <= pause_getI3574;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1546_forever6893377\;
            end case;
          when pause_getII3585 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1494\ := \$arr3399_value\;
            \$v3583\ := \$arr3400_ptr_take\;
            if \$v3583\(0) = '1' then
              \state\ <= q_wait3582;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3580;
            end if;
          when pause_getII3589 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1551\ := \$arr3400_value\;
            \$v3587\ := \$arr3399_ptr_take\;
            if \$v3587\(0) = '1' then
              \state\ <= q_wait3586;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1551\));
              \state\ <= pause_getI3584;
            end if;
          when pause_getII3602 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3302\ := \$arr3399_value\;
            eclat_print_string(of_string("[ "));
            
            \$1371_show_rib6323365_arg\ := \$v3302\(0 to 35) & \$1371_show_rib6323365_arg\(36 to 67) & eclat_add(\$1371_show_rib6323365_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$1371_show_rib6323365\;
          when pause_getII3611 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1394\ := \$arr3400_value\;
            \$1393\ := "0010" & \$1394\;
            \$1370\ := \$1393\ & "00000000000000000000000000000011" & "00000000000000000000000000000000";
            \$1371_show_rib6323365_arg\ := \$1370\;
            \state\ <= \$1371_show_rib6323365\;
          when pause_getII3630 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2916\ := \$arr3399_value\;
            \$1405\ := \$v2916\(72 to 107);
            \$v3626\ := \$1405\;
            \$v3627\ := \$v3626\(0 to 3);
            \$v3625\ := \$v3626\(4 to 35);
            case \$v3627\ is
            when "0010" =>
              \$1406_i\ := \$v3625\(0 to 31);
              \$1404\ := \$1406_i\;
              \$v3624\ := \$arr3401_ptr_take\;
              if \$v3624\(0) = '1' then
                \state\ <= q_wait3623;
              else
                \$arr3401_ptr_take\(0) := '1';
                \$arr3401_ptr_write\ <= 0;
                \$arr3401_write_request\ <= '1';
                \$arr3401_write\ <= \$1404\;
                \state\ <= pause_setI3621;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1410_forever6893367\;
            end case;
          when pause_getII3638 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3315\ := \$arr3399_value\;
            eclat_print_string(of_string("["));
            
            \$1423_print_value6133369_arg\ := \$v3315\(0 to 35);
            \state\ <= \$1423_print_value6133369\;
          when pause_getII3647 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2920\ := \$arr3399_value\;
            \$1422\ := \$v2920\(72 to 107);
            \$1423_print_value6133369_arg\ := \$1422\;
            \state\ <= \$1423_print_value6133369\;
          when pause_getII3657 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1492\ := \$arr3400_value\;
            \$1491\ := "0010" & \$1492\;
            \$1490\ := \$1491\ & \$1486\(36 to 71) & \$1073_loop667_arg\(68 to 103);
            \$v3655\ := \$arr3399_ptr_take\;
            if \$v3655\(0) = '1' then
              \state\ <= q_wait3654;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1490\;
              \state\ <= pause_setI3652;
            end if;
          when pause_getII3661 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1486\ := \$arr3399_value\;
            \$v3659\ := \$arr3400_ptr_take\;
            if \$v3659\(0) = '1' then
              \state\ <= q_wait3658;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3656;
            end if;
          when pause_getII3670 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2925\ := \$arr3399_value\;
            \$1445\ := \$v2925\(72 to 107);
            \$1443\ := \$1444\ & \$1439\(36 to 71) & \$1445\;
            \$v3667\ := \$arr3399_ptr_take\;
            if \$v3667\(0) = '1' then
              \state\ <= q_wait3666;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1443\;
              \state\ <= pause_setI3664;
            end if;
          when pause_getII3677 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2929\ := \$arr3399_value\;
            \$1444\ := \$v2929\(0 to 35);
            \$v3673\ := \$1438_k\;
            \$v3674\ := \$v3673\(0 to 3);
            \$v3668\ := \$v3673\(4 to 35);
            case \$v3674\ is
            when "0010" =>
              \$1446_t\ := \$v3668\(0 to 31);
              \$v3672\ := \$arr3399_ptr_take\;
              if \$v3672\(0) = '1' then
                \state\ <= q_wait3671;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1446_t\));
                \state\ <= pause_getI3669;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1450_forever6893371\;
            end case;
          when pause_getII3683 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1439\ := \$arr3399_value\;
            \$v3680\ := \$1438_k\;
            \$v3681\ := \$v3680\(0 to 3);
            \$v3675\ := \$v3680\(4 to 35);
            case \$v3681\ is
            when "0010" =>
              \$1454_t\ := \$v3675\(0 to 31);
              \$v3679\ := \$arr3399_ptr_take\;
              if \$v3679\(0) = '1' then
                \state\ <= q_wait3678;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1454_t\));
                \state\ <= pause_getI3676;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1458_forever6893372\;
            end case;
          when pause_getII3697 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3302\ := \$arr3399_value\;
            eclat_print_string(of_string("[ "));
            
            \$411_show_rib6323357_arg\ := \$v3302\(0 to 35) & \$411_show_rib6323357_arg\(36 to 67) & eclat_add(\$411_show_rib6323357_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$411_show_rib6323357\;
          when pause_getII3707 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2985\ := \$arr3399_value\;
            \$v402\ := \$v2985\(36 to 71);
            \$1464_loop6693373_arg\ := \$v402\;
            \state\ <= \$1464_loop6693373\;
          when pause_getII3722 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3302\ := \$arr3399_value\;
            eclat_print_string(of_string("[ "));
            
            \$411_show_rib6323359_arg\ := \$v3302\(0 to 35) & \$411_show_rib6323359_arg\(36 to 67) & eclat_add(\$411_show_rib6323359_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$411_show_rib6323359\;
          when pause_getII3734 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v2989\ := \$arr3399_value\;
            \$1467_tag\ := \$v2989\(72 to 107);
            \$v3730\ := \$1467_tag\;
            \$v3731\ := \$v3730\(0 to 3);
            \$v3686\ := \$v3730\(4 to 35);
            case \$v3731\ is
            when "0010" =>
              \$411_show_rib6323357_arg\ := \$1464_loop6693373_arg\ & "00000000000000000000000000000101" & "00000000000000000000000000000000";
              \state\ <= \$411_show_rib6323357\;
            when "0001" =>
              \$411_show_rib6323359_arg\ := \$1464_loop6693373_arg\ & "00000000000000000000000000000101" & "00000000000000000000000000000000";
              \state\ <= \$411_show_rib6323359\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cont 2"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1473_forever6893356\;
            end case;
          when pause_getII3740 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1485\ := \$arr3400_value\;
            \$1463\ := "0010" & \$1485\;
            \$1464_loop6693373_arg\ := \$1463\;
            \state\ <= \$1464_loop6693373\;
          when pause_getII3757 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1656\ := \$arr3399_value\;
            \$1108\ := \$v1656\(36 to 71);
            \$v3753\ := \$1108\;
            \$v3754\ := \$v3753\(0 to 3);
            \$v3752\ := \$v3753\(4 to 35);
            case \$v3754\ is
            when "0010" =>
              \$1109_i\ := \$v3752\(0 to 31);
              \$1107\ := \$1109_i\;
              \$v3751\ := \$arr3402_ptr_take\;
              if \$v3751\(0) = '1' then
                \state\ <= q_wait3750;
              else
                \$arr3402_ptr_take\(0) := '1';
                \$arr3402_ptr_write\ <= 0;
                \$arr3402_write_request\ <= '1';
                \$arr3402_write\ <= \$1107\;
                \state\ <= pause_setI3748;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1113_forever6893378\;
            end case;
          when pause_getII3763 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1126\ := \$arr3402_value\;
            \$1117\ := "0010" & \$1126\;
            \$v3760\ := \$1117\;
            \$v3761\ := \$v3760\(0 to 3);
            \$v3755\ := \$v3760\(4 to 35);
            case \$v3761\ is
            when "0010" =>
              \$1118_t\ := \$v3755\(0 to 31);
              \$v3759\ := \$arr3399_ptr_take\;
              if \$v3759\(0) = '1' then
                \state\ <= q_wait3758;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1118_t\));
                \state\ <= pause_getI3756;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1122_forever6893379\;
            end case;
          when pause_getII3775 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1102\ := \$arr3399_value\;
            \$v3772\ := \$1101_car\;
            \$v3773\ := \$v3772\(0 to 3);
            \$v3771\ := \$v3772\(4 to 35);
            case \$v3773\ is
            when "0010" =>
              \$1130_i\ := \$v3771\(0 to 31);
              \$1127\ := \$1130_i\;
              \$v3770\ := \$arr3399_ptr_take\;
              if \$v3770\(0) = '1' then
                \state\ <= q_wait3769;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$v3766\ := "00000000000000000000000000000010";
                \$arr3399_ptr_write\ <= to_integer(unsigned(\$1127\));
                \$arr3399_write_request\ <= '1';
                \$arr3399_write\ <= "0010" & \$v3766\ & \$1102\(36 to 71) & \$1102\(72 to 107);
                \state\ <= pause_setI3767;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1134_forever6893380\;
            end case;
          when pause_getII3783 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1666\ := \$arr3399_value\;
            \$1101_car\ := \$v1666\(0 to 35);
            \$v3779\ := \$1101_car\;
            \$v3780\ := \$v3779\(0 to 3);
            \$v3778\ := \$v3779\(4 to 35);
            case \$v3780\ is
            when "0010" =>
              \$1139_i\ := \$v3778\(0 to 31);
              \$1138\ := \$1139_i\;
              \$v3777\ := \$arr3399_ptr_take\;
              if \$v3777\(0) = '1' then
                \state\ <= q_wait3776;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1138\));
                \state\ <= pause_getI3774;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1143_forever6893381\;
            end case;
          when pause_getII3789 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1156\ := \$arr3402_value\;
            \$1147\ := "0010" & \$1156\;
            \$v3786\ := \$1147\;
            \$v3787\ := \$v3786\(0 to 3);
            \$v3781\ := \$v3786\(4 to 35);
            case \$v3787\ is
            when "0010" =>
              \$1148_t\ := \$v3781\(0 to 31);
              \$v3785\ := \$arr3399_ptr_take\;
              if \$v3785\(0) = '1' then
                \state\ <= q_wait3784;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1148_t\));
                \state\ <= pause_getI3782;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1152_forever6893382\;
            end case;
          when pause_getII3801 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1675\ := \$arr3399_value\;
            \$1164\ := \$v1675\(36 to 71);
            \$v3797\ := \$1164\;
            \$v3798\ := \$v3797\(0 to 3);
            \$v3796\ := \$v3797\(4 to 35);
            case \$v3798\ is
            when "0010" =>
              \$1165_i\ := \$v3796\(0 to 31);
              \$1163\ := \$1165_i\;
              \$v3795\ := \$arr3402_ptr_take\;
              if \$v3795\(0) = '1' then
                \state\ <= q_wait3794;
              else
                \$arr3402_ptr_take\(0) := '1';
                \$arr3402_ptr_write\ <= 0;
                \$arr3402_write_request\ <= '1';
                \$arr3402_write\ <= \$1163\;
                \state\ <= pause_setI3792;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1169_forever6893383\;
            end case;
          when pause_getII3807 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1182\ := \$arr3402_value\;
            \$1173\ := "0010" & \$1182\;
            \$v3804\ := \$1173\;
            \$v3805\ := \$v3804\(0 to 3);
            \$v3799\ := \$v3804\(4 to 35);
            case \$v3805\ is
            when "0010" =>
              \$1174_t\ := \$v3799\(0 to 31);
              \$v3803\ := \$arr3399_ptr_take\;
              if \$v3803\(0) = '1' then
                \state\ <= q_wait3802;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1174_t\));
                \state\ <= pause_getI3800;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1178_forever6893384\;
            end case;
          when pause_getII3819 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1158\ := \$arr3399_value\;
            \$v3816\ := \$1157_car\;
            \$v3817\ := \$v3816\(0 to 3);
            \$v3815\ := \$v3816\(4 to 35);
            case \$v3817\ is
            when "0010" =>
              \$1186_i\ := \$v3815\(0 to 31);
              \$1183\ := \$1186_i\;
              \$v3814\ := \$arr3399_ptr_take\;
              if \$v3814\(0) = '1' then
                \state\ <= q_wait3813;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$v3810\ := "00000000000000000000000000000001";
                \$arr3399_ptr_write\ <= to_integer(unsigned(\$1183\));
                \$arr3399_write_request\ <= '1';
                \$arr3399_write\ <= "0010" & \$v3810\ & \$1158\(36 to 71) & \$1158\(72 to 107);
                \state\ <= pause_setI3811;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1190_forever6893385\;
            end case;
          when pause_getII3827 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1685\ := \$arr3399_value\;
            \$1157_car\ := \$v1685\(0 to 35);
            \$v3823\ := \$1157_car\;
            \$v3824\ := \$v3823\(0 to 3);
            \$v3822\ := \$v3823\(4 to 35);
            case \$v3824\ is
            when "0010" =>
              \$1195_i\ := \$v3822\(0 to 31);
              \$1194\ := \$1195_i\;
              \$v3821\ := \$arr3399_ptr_take\;
              if \$v3821\(0) = '1' then
                \state\ <= q_wait3820;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1194\));
                \state\ <= pause_getI3818;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1199_forever6893386\;
            end case;
          when pause_getII3833 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1212\ := \$arr3402_value\;
            \$1203\ := "0010" & \$1212\;
            \$v3830\ := \$1203\;
            \$v3831\ := \$v3830\(0 to 3);
            \$v3825\ := \$v3830\(4 to 35);
            case \$v3831\ is
            when "0010" =>
              \$1204_t\ := \$v3825\(0 to 31);
              \$v3829\ := \$arr3399_ptr_take\;
              if \$v3829\(0) = '1' then
                \state\ <= q_wait3828;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1204_t\));
                \state\ <= pause_getI3826;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1208_forever6893387\;
            end case;
          when pause_getII3845 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1694\ := \$arr3399_value\;
            \$1220\ := \$v1694\(36 to 71);
            \$v3841\ := \$1220\;
            \$v3842\ := \$v3841\(0 to 3);
            \$v3840\ := \$v3841\(4 to 35);
            case \$v3842\ is
            when "0010" =>
              \$1221_i\ := \$v3840\(0 to 31);
              \$1219\ := \$1221_i\;
              \$v3839\ := \$arr3402_ptr_take\;
              if \$v3839\(0) = '1' then
                \state\ <= q_wait3838;
              else
                \$arr3402_ptr_take\(0) := '1';
                \$arr3402_ptr_write\ <= 0;
                \$arr3402_write_request\ <= '1';
                \$arr3402_write\ <= \$1219\;
                \state\ <= pause_setI3836;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1225_forever6893388\;
            end case;
          when pause_getII3851 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1238\ := \$arr3402_value\;
            \$1229\ := "0010" & \$1238\;
            \$v3848\ := \$1229\;
            \$v3849\ := \$v3848\(0 to 3);
            \$v3843\ := \$v3848\(4 to 35);
            case \$v3849\ is
            when "0010" =>
              \$1230_t\ := \$v3843\(0 to 31);
              \$v3847\ := \$arr3399_ptr_take\;
              if \$v3847\(0) = '1' then
                \state\ <= q_wait3846;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1230_t\));
                \state\ <= pause_getI3844;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1234_forever6893389\;
            end case;
          when pause_getII3863 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1214\ := \$arr3399_value\;
            \$v3860\ := \$1213_car\;
            \$v3861\ := \$v3860\(0 to 3);
            \$v3859\ := \$v3860\(4 to 35);
            case \$v3861\ is
            when "0010" =>
              \$1242_i\ := \$v3859\(0 to 31);
              \$1239\ := \$1242_i\;
              \$v3858\ := \$arr3399_ptr_take\;
              if \$v3858\(0) = '1' then
                \state\ <= q_wait3857;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$v3854\ := "00000000000000000000000000000011";
                \$arr3399_ptr_write\ <= to_integer(unsigned(\$1239\));
                \$arr3399_write_request\ <= '1';
                \$arr3399_write\ <= "0010" & \$v3854\ & \$1214\(36 to 71) & \$1214\(72 to 107);
                \state\ <= pause_setI3855;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1246_forever6893390\;
            end case;
          when pause_getII3871 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1704\ := \$arr3399_value\;
            \$1213_car\ := \$v1704\(0 to 35);
            \$v3867\ := \$1213_car\;
            \$v3868\ := \$v3867\(0 to 3);
            \$v3866\ := \$v3867\(4 to 35);
            case \$v3868\ is
            when "0010" =>
              \$1251_i\ := \$v3866\(0 to 31);
              \$1250\ := \$1251_i\;
              \$v3865\ := \$arr3399_ptr_take\;
              if \$v3865\(0) = '1' then
                \state\ <= q_wait3864;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1250\));
                \state\ <= pause_getI3862;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1255_forever6893391\;
            end case;
          when pause_getII3877 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1268\ := \$arr3402_value\;
            \$1259\ := "0010" & \$1268\;
            \$v3874\ := \$1259\;
            \$v3875\ := \$v3874\(0 to 3);
            \$v3869\ := \$v3874\(4 to 35);
            case \$v3875\ is
            when "0010" =>
              \$1260_t\ := \$v3869\(0 to 31);
              \$v3873\ := \$arr3399_ptr_take\;
              if \$v3873\(0) = '1' then
                \state\ <= q_wait3872;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1260_t\));
                \state\ <= pause_getI3870;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1264_forever6893392\;
            end case;
          when pause_getII3889 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1713\ := \$arr3399_value\;
            \$1276\ := \$v1713\(36 to 71);
            \$v3885\ := \$1276\;
            \$v3886\ := \$v3885\(0 to 3);
            \$v3884\ := \$v3885\(4 to 35);
            case \$v3886\ is
            when "0010" =>
              \$1277_i\ := \$v3884\(0 to 31);
              \$1275\ := \$1277_i\;
              \$v3883\ := \$arr3402_ptr_take\;
              if \$v3883\(0) = '1' then
                \state\ <= q_wait3882;
              else
                \$arr3402_ptr_take\(0) := '1';
                \$arr3402_ptr_write\ <= 0;
                \$arr3402_write_request\ <= '1';
                \$arr3402_write\ <= \$1275\;
                \state\ <= pause_setI3880;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1281_forever6893393\;
            end case;
          when pause_getII3895 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1294\ := \$arr3402_value\;
            \$1285\ := "0010" & \$1294\;
            \$v3892\ := \$1285\;
            \$v3893\ := \$v3892\(0 to 3);
            \$v3887\ := \$v3892\(4 to 35);
            case \$v3893\ is
            when "0010" =>
              \$1286_t\ := \$v3887\(0 to 31);
              \$v3891\ := \$arr3399_ptr_take\;
              if \$v3891\(0) = '1' then
                \state\ <= q_wait3890;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1286_t\));
                \state\ <= pause_getI3888;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1290_forever6893394\;
            end case;
          when pause_getII3907 =>
            \$arr3399_ptr_take\(0) := '0';
            \$1270\ := \$arr3399_value\;
            \$v3904\ := \$1269_car\;
            \$v3905\ := \$v3904\(0 to 3);
            \$v3903\ := \$v3904\(4 to 35);
            case \$v3905\ is
            when "0010" =>
              \$1298_i\ := \$v3903\(0 to 31);
              \$1295\ := \$1298_i\;
              \$v3902\ := \$arr3399_ptr_take\;
              if \$v3902\(0) = '1' then
                \state\ <= q_wait3901;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$v3898\ := "00000000000000000000000000000000";
                \$arr3399_ptr_write\ <= to_integer(unsigned(\$1295\));
                \$arr3399_write_request\ <= '1';
                \$arr3399_write\ <= "0010" & \$v3898\ & \$1270\(36 to 71) & \$1270\(72 to 107);
                \state\ <= pause_setI3899;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1302_forever6893395\;
            end case;
          when pause_getII3915 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v1723\ := \$arr3399_value\;
            \$1269_car\ := \$v1723\(0 to 35);
            \$v3911\ := \$1269_car\;
            \$v3912\ := \$v3911\(0 to 3);
            \$v3910\ := \$v3911\(4 to 35);
            case \$v3912\ is
            when "0010" =>
              \$1307_i\ := \$v3910\(0 to 31);
              \$1306\ := \$1307_i\;
              \$v3909\ := \$arr3399_ptr_take\;
              if \$v3909\(0) = '1' then
                \state\ <= q_wait3908;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1306\));
                \state\ <= pause_getI3906;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1311_forever6893396\;
            end case;
          when pause_getII3921 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1324\ := \$arr3402_value\;
            \$1315\ := "0010" & \$1324\;
            \$v3918\ := \$1315\;
            \$v3919\ := \$v3918\(0 to 3);
            \$v3913\ := \$v3918\(4 to 35);
            case \$v3919\ is
            when "0010" =>
              \$1316_t\ := \$v3913\(0 to 31);
              \$v3917\ := \$arr3399_ptr_take\;
              if \$v3917\(0) = '1' then
                \state\ <= q_wait3916;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1316_t\));
                \state\ <= pause_getI3914;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1320_forever6893397\;
            end case;
          when pause_getII3929 =>
            \$arr3400_ptr_take\(0) := '0';
            \$1325\ := \$arr3400_value\;
            \$v3927\ := \$arr3404_ptr_take\;
            if \$v3927\(0) = '1' then
              \state\ <= q_wait3926;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= \$1325\;
              \state\ <= pause_setI3924;
            end if;
          when pause_getII3937 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1326\ := \$arr3402_value\;
            \$v3935\ := \$arr3401_ptr_take\;
            if \$v3935\(0) = '1' then
              \state\ <= q_wait3934;
            else
              \$arr3401_ptr_take\(0) := '1';
              \$arr3401_ptr_write\ <= 0;
              \$arr3401_write_request\ <= '1';
              \$arr3401_write\ <= \$1326\;
              \state\ <= pause_setI3932;
            end if;
          when pause_getII3947 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1336\ := \$arr3402_value\;
            \$1333\ := "0010" & \$1336\;
            \$v3944\ := "00000000000000000000000000000000";
            \$v3945\ := "00000000000000000000000000000001";
            \$1328\ := "0001" & \$v3944\ & \$1333\ & "0001" & \$v3945\;
            \$1327\ := \$1328\(0 to 35) & \$1328\(36 to 71) & \$1328\(72 to 107);
            \$v3943\ := \$arr3399_ptr_take\;
            if \$v3943\(0) = '1' then
              \state\ <= q_wait3942;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= 0;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1327\;
              \state\ <= pause_setI3940;
            end if;
          when pause_getII3955 =>
            \$arr3402_ptr_take\(0) := '0';
            \$1337\ := \$arr3402_value\;
            \$v3953\ := \$arr3404_ptr_take\;
            if \$v3953\(0) = '1' then
              \state\ <= q_wait3952;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= \$1337\;
              \state\ <= pause_setI3950;
            end if;
          when pause_setI3427 =>
            \$arr3403_write_request\ <= '0';
            \state\ <= pause_setII3428;
          when pause_setI3447 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII3448;
          when pause_setI3452 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3453;
          when pause_setI3460 =>
            \$arr3400_write_request\ <= '0';
            \state\ <= pause_setII3461;
          when pause_setI3504 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3505;
          when pause_setI3508 =>
            \$arr3400_write_request\ <= '0';
            \state\ <= pause_setII3509;
          when pause_setI3516 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII3517;
          when pause_setI3520 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3521;
          when pause_setI3538 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII3539;
          when pause_setI3543 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3544;
          when pause_setI3551 =>
            \$arr3400_write_request\ <= '0';
            \state\ <= pause_setII3552;
          when pause_setI3614 =>
            \$arr3400_write_request\ <= '0';
            \state\ <= pause_setII3615;
          when pause_setI3621 =>
            \$arr3401_write_request\ <= '0';
            \state\ <= pause_setII3622;
          when pause_setI3652 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3653;
          when pause_setI3664 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3665;
          when pause_setI3748 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII3749;
          when pause_setI3767 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3768;
          when pause_setI3792 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII3793;
          when pause_setI3811 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3812;
          when pause_setI3836 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII3837;
          when pause_setI3855 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3856;
          when pause_setI3880 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII3881;
          when pause_setI3899 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3900;
          when pause_setI3924 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII3925;
          when pause_setI3932 =>
            \$arr3401_write_request\ <= '0';
            \state\ <= pause_setII3933;
          when pause_setI3940 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3941;
          when pause_setI3950 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII3951;
          when pause_setI3958 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII3959;
          when pause_setI3965 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3966;
          when pause_setI3972 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3973;
          when pause_setI3979 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3980;
          when pause_setI3986 =>
            \$arr3399_write_request\ <= '0';
            \state\ <= pause_setII3987;
          when pause_setI3990 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII3991;
          when pause_setI3994 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII3995;
          when pause_setI3998 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII3999;
          when pause_setI4002 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII4003;
          when pause_setI4006 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII4007;
          when pause_setI4010 =>
            \$arr3405_write_request\ <= '0';
            \state\ <= pause_setII4011;
          when pause_setI4014 =>
            \$arr3404_write_request\ <= '0';
            \state\ <= pause_setII4015;
          when pause_setI4018 =>
            \$arr3403_write_request\ <= '0';
            \state\ <= pause_setII4019;
          when pause_setI4022 =>
            \$arr3402_write_request\ <= '0';
            \state\ <= pause_setII4023;
          when pause_setI4026 =>
            \$arr3400_write_request\ <= '0';
            \state\ <= pause_setII4027;
          when pause_setI4030 =>
            \$arr3401_write_request\ <= '0';
            \state\ <= pause_setII4031;
          when pause_setII3428 =>
            \$arr3403_ptr_take\(0) := '0';
            \$1651\ := \$1653_c\;
            \$1650\ := \$1651\ & X"000000" & X"23";
            \$1648_x\ := eclat_sub(\$1650\);
            \$1638_x\ := eclat_if(eclat_lt(\$1648_x\ & "00000000000000000000000000000000") & X"000000" & X"39" & \$1648_x\);
            \$v3426\ := eclat_lt(\$1638_x\ & X"000000" & X"2e");
            if \$v3426\(0) = '1' then
              \state\ <= \$1070_get_int640\;
            else
              \$1070_get_int640_arg\ := eclat_sub(eclat_add(eclat_mult(\$1070_get_int640_arg\ & X"000000" & X"2e") & \$1638_x\) & X"000000" & X"2e");
              \state\ <= \$1070_get_int640\;
            end if;
          when pause_setII3448 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v3446\ := \$arr3404_ptr_take\;
            if \$v3446\(0) = '1' then
              \state\ <= q_wait3445;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3443;
            end if;
          when pause_setII3453 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3450\ := \$arr3404_ptr_take\;
            if \$v3450\(0) = '1' then
              \state\ <= q_wait3449;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1588_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3447;
            end if;
          when pause_setII3461 =>
            \$arr3400_ptr_take\(0) := '0';
            \$v3459\ := \$arr3404_ptr_take\;
            if \$v3459\(0) = '1' then
              \state\ <= q_wait3458;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3456;
            end if;
          when pause_setII3505 =>
            \$arr3399_ptr_take\(0) := '0';
            \state\ <= \$1072_rest_loop668\;
          when pause_setII3509 =>
            \$arr3400_ptr_take\(0) := '0';
            \$v3507\ := \$arr3399_ptr_take\;
            if \$v3507\(0) = '1' then
              \state\ <= q_wait3506;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3501\ := eclat_add(\$1072_rest_loop668_arg\(100 to 131) & "00000000000000000000000000000001");
              \$v3502\ := "00000000000000000000000000000000";
              \$v3503\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1072_rest_loop668_arg\(68 to 99)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3501\ & "0001" & \$v3502\ & "0001" & \$v3503\;
              \state\ <= pause_setI3504;
            end if;
          when pause_setII3517 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v3515\ := \$arr3404_ptr_take\;
            if \$v3515\(0) = '1' then
              \state\ <= q_wait3514;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3512;
            end if;
          when pause_setII3521 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3519\ := \$arr3404_ptr_take\;
            if \$v3519\(0) = '1' then
              \state\ <= q_wait3518;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1571_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3516;
            end if;
          when pause_setII3539 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v3537\ := \$arr3404_ptr_take\;
            if \$v3537\(0) = '1' then
              \state\ <= q_wait3536;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3534;
            end if;
          when pause_setII3544 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3541\ := \$arr3404_ptr_take\;
            if \$v3541\(0) = '1' then
              \state\ <= q_wait3540;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1504_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3538;
            end if;
          when pause_setII3552 =>
            \$arr3400_ptr_take\(0) := '0';
            \$v3550\ := \$arr3404_ptr_take\;
            if \$v3550\(0) = '1' then
              \state\ <= q_wait3549;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3547;
            end if;
          when pause_setII3615 =>
            \$arr3400_ptr_take\(0) := '0';
            \$v3613\ := \$arr3400_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3610;
            end if;
          when pause_setII3622 =>
            \$arr3401_ptr_take\(0) := '0';
            \$v3619\ := \$1073_loop667_arg\(32 to 67);
            \$v3620\ := \$v3619\(0 to 3);
            \$v3618\ := \$v3619\(4 to 35);
            case \$v3620\ is
            when "0010" =>
              \$1396_i\ := \$v3618\(0 to 31);
              \$1395\ := \$1396_i\;
              \$v3617\ := \$arr3400_ptr_take\;
              if \$v3617\(0) = '1' then
                \state\ <= q_wait3616;
              else
                \$arr3400_ptr_take\(0) := '1';
                \$arr3400_ptr_write\ <= 0;
                \$arr3400_write_request\ <= '1';
                \$arr3400_write\ <= \$1395\;
                \state\ <= pause_setI3614;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1400_forever6893366\;
            end case;
          when pause_setII3653 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3650\ := \$1073_loop667_arg\(104 to 139);
            \$v3651\ := \$v3650\(0 to 3);
            \$v3645\ := \$v3650\(4 to 35);
            case \$v3651\ is
            when "0010" =>
              \$1429_t\ := \$v3645\(0 to 31);
              \$v3649\ := \$arr3399_ptr_take\;
              if \$v3649\(0) = '1' then
                \state\ <= q_wait3648;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1429_t\));
                \state\ <= pause_getI3646;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1433_forever6893370\;
            end case;
          when pause_setII3665 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3650\ := \$1073_loop667_arg\(104 to 139);
            \$v3651\ := \$v3650\(0 to 3);
            \$v3645\ := \$v3650\(4 to 35);
            case \$v3651\ is
            when "0010" =>
              \$1429_t\ := \$v3645\(0 to 31);
              \$v3649\ := \$arr3399_ptr_take\;
              if \$v3649\(0) = '1' then
                \state\ <= q_wait3648;
              else
                \$arr3399_ptr_take\(0) := '1';
                \$arr3399_ptr\ <= to_integer(unsigned(\$1429_t\));
                \state\ <= pause_getI3646;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1433_forever6893370\;
            end case;
          when pause_setII3749 =>
            \$arr3402_ptr_take\(0) := '0';
            eclat_print_string(of_string("Compilation reussi, pas de bug dans la syntaxe "));
            
            result3406 := eclat_unit;
            eclat_print_newline(eclat_unit);
            
            rdy3407 := eclat_true;
            \state\ <= compute3408;
          when pause_setII3768 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3765\ := \$arr3402_ptr_take\;
            if \$v3765\(0) = '1' then
              \state\ <= q_wait3764;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3762;
            end if;
          when pause_setII3793 =>
            \$arr3402_ptr_take\(0) := '0';
            \$v3791\ := \$arr3402_ptr_take\;
            if \$v3791\(0) = '1' then
              \state\ <= q_wait3790;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3788;
            end if;
          when pause_setII3812 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3809\ := \$arr3402_ptr_take\;
            if \$v3809\(0) = '1' then
              \state\ <= q_wait3808;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3806;
            end if;
          when pause_setII3837 =>
            \$arr3402_ptr_take\(0) := '0';
            \$v3835\ := \$arr3402_ptr_take\;
            if \$v3835\(0) = '1' then
              \state\ <= q_wait3834;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3832;
            end if;
          when pause_setII3856 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3853\ := \$arr3402_ptr_take\;
            if \$v3853\(0) = '1' then
              \state\ <= q_wait3852;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3850;
            end if;
          when pause_setII3881 =>
            \$arr3402_ptr_take\(0) := '0';
            \$v3879\ := \$arr3402_ptr_take\;
            if \$v3879\(0) = '1' then
              \state\ <= q_wait3878;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3876;
            end if;
          when pause_setII3900 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3897\ := \$arr3402_ptr_take\;
            if \$v3897\(0) = '1' then
              \state\ <= q_wait3896;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3894;
            end if;
          when pause_setII3925 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v3923\ := \$arr3402_ptr_take\;
            if \$v3923\(0) = '1' then
              \state\ <= q_wait3922;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3920;
            end if;
          when pause_setII3933 =>
            \$arr3401_ptr_take\(0) := '0';
            \$v3931\ := \$arr3400_ptr_take\;
            if \$v3931\(0) = '1' then
              \state\ <= q_wait3930;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3928;
            end if;
          when pause_setII3941 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3939\ := \$arr3402_ptr_take\;
            if \$v3939\(0) = '1' then
              \state\ <= q_wait3938;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3936;
            end if;
          when pause_setII3951 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v3949\ := \$arr3402_ptr_take\;
            if \$v3949\(0) = '1' then
              \state\ <= q_wait3948;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3946;
            end if;
          when pause_setII3959 =>
            \$arr3402_ptr_take\(0) := '0';
            \$v3957\ := \$arr3402_ptr_take\;
            if \$v3957\(0) = '1' then
              \state\ <= q_wait3956;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3954;
            end if;
          when pause_setII3966 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3961\ := \$arr3402_ptr_take\;
            if \$v3961\(0) = '1' then
              \state\ <= q_wait3960;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= "00000000000000000000000000000011";
              \state\ <= pause_setI3958;
            end if;
          when pause_setII3973 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3968\ := \$arr3399_ptr_take\;
            if \$v3968\(0) = '1' then
              \state\ <= q_wait3967;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3962\ := "00000000000000000000000000000001";
              \$v3963\ := "00000000000000000000000000000010";
              \$v3964\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 3;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3962\ & "0010" & \$v3963\ & "0001" & \$v3964\;
              \state\ <= pause_setI3965;
            end if;
          when pause_setII3980 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3975\ := \$arr3399_ptr_take\;
            if \$v3975\(0) = '1' then
              \state\ <= q_wait3974;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3969\ := "00000000000000000000000000000000";
              \$v3970\ := "00000000000000000000000000000000";
              \$v3971\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 2;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3969\ & "0001" & \$v3970\ & "0001" & \$v3971\;
              \state\ <= pause_setI3972;
            end if;
          when pause_setII3987 =>
            \$arr3399_ptr_take\(0) := '0';
            \$v3982\ := \$arr3399_ptr_take\;
            if \$v3982\(0) = '1' then
              \state\ <= q_wait3981;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3976\ := "00000000000000000000000000000000";
              \$v3977\ := "00000000000000000000000000000000";
              \$v3978\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 1;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3976\ & "0001" & \$v3977\ & "0001" & \$v3978\;
              \state\ <= pause_setI3979;
            end if;
          when pause_setII3991 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v3989\ := \$arr3399_ptr_take\;
            if \$v3989\(0) = '1' then
              \state\ <= q_wait3988;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3983\ := "00000000000000000000000000000000";
              \$v3984\ := "00000000000000000000000000000000";
              \$v3985\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 0;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3983\ & "0001" & \$v3984\ & "0001" & \$v3985\;
              \state\ <= pause_setI3986;
            end if;
          when pause_setII3995 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v3993\ := \$arr3405_ptr_take\;
            if \$v3993\(0) = '1' then
              \state\ <= q_wait3992;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 5;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI3990;
            end if;
          when pause_setII3999 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v3997\ := \$arr3405_ptr_take\;
            if \$v3997\(0) = '1' then
              \state\ <= q_wait3996;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 4;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI3994;
            end if;
          when pause_setII4003 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v4001\ := \$arr3405_ptr_take\;
            if \$v4001\(0) = '1' then
              \state\ <= q_wait4000;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 3;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI3998;
            end if;
          when pause_setII4007 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v4005\ := \$arr3405_ptr_take\;
            if \$v4005\(0) = '1' then
              \state\ <= q_wait4004;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 2;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4002;
            end if;
          when pause_setII4011 =>
            \$arr3405_ptr_take\(0) := '0';
            \$v4009\ := \$arr3405_ptr_take\;
            if \$v4009\(0) = '1' then
              \state\ <= q_wait4008;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 1;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI4006;
            end if;
          when pause_setII4015 =>
            \$arr3404_ptr_take\(0) := '0';
            \$v4013\ := \$arr3405_ptr_take\;
            if \$v4013\(0) = '1' then
              \state\ <= q_wait4012;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 0;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= X"000000" & X"14";
              \state\ <= pause_setI4010;
            end if;
          when pause_setII4019 =>
            \$arr3403_ptr_take\(0) := '0';
            \$v4017\ := \$arr3404_ptr_take\;
            if \$v4017\(0) = '1' then
              \state\ <= q_wait4016;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4014;
            end if;
          when pause_setII4023 =>
            \$arr3402_ptr_take\(0) := '0';
            \$v4021\ := \$arr3403_ptr_take\;
            if \$v4021\(0) = '1' then
              \state\ <= q_wait4020;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr_write\ <= 0;
              \$arr3403_write_request\ <= '1';
              \$arr3403_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4018;
            end if;
          when pause_setII4027 =>
            \$arr3400_ptr_take\(0) := '0';
            \$v4025\ := \$arr3402_ptr_take\;
            if \$v4025\(0) = '1' then
              \state\ <= q_wait4024;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4022;
            end if;
          when pause_setII4031 =>
            \$arr3401_ptr_take\(0) := '0';
            \$v4029\ := \$arr3400_ptr_take\;
            if \$v4029\(0) = '1' then
              \state\ <= q_wait4028;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI4026;
            end if;
          when q_wait3415 =>
            \$v3416\ := \$arr3399_ptr_take\;
            if \$v3416\(0) = '1' then
              \state\ <= q_wait3415;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1069_list_tail637_arg\(0 to 31)));
              \state\ <= pause_getI3413;
            end if;
          when q_wait3423 =>
            \$v3424\ := \$arr3399_ptr_take\;
            if \$v3424\(0) = '1' then
              \state\ <= q_wait3423;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1069_list_tail637_arg\(0 to 31)));
              \state\ <= pause_getI3421;
            end if;
          when q_wait3429 =>
            \$v3430\ := \$arr3403_ptr_take\;
            if \$v3430\(0) = '1' then
              \state\ <= q_wait3429;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr_write\ <= 0;
              \$arr3403_write_request\ <= '1';
              \$arr3403_write\ <= \$1655\;
              \state\ <= pause_setI3427;
            end if;
          when q_wait3433 =>
            \$v3434\ := \$arr3403_ptr_take\;
            if \$v3434\(0) = '1' then
              \state\ <= q_wait3433;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr\ <= 0;
              \state\ <= pause_getI3431;
            end if;
          when q_wait3437 =>
            \$v3438\ := \$arr3398_ptr_take\;
            if \$v3438\(0) = '1' then
              \state\ <= q_wait3437;
            else
              \$arr3398_ptr_take\(0) := '1';
              \$arr3398_ptr\ <= to_integer(unsigned(\$1658\));
              \state\ <= pause_getI3435;
            end if;
          when q_wait3441 =>
            \$v3442\ := \$arr3403_ptr_take\;
            if \$v3442\(0) = '1' then
              \state\ <= q_wait3441;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr\ <= 0;
              \state\ <= pause_getI3439;
            end if;
          when q_wait3445 =>
            \$v3446\ := \$arr3404_ptr_take\;
            if \$v3446\(0) = '1' then
              \state\ <= q_wait3445;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3443;
            end if;
          when q_wait3449 =>
            \$v3450\ := \$arr3404_ptr_take\;
            if \$v3450\(0) = '1' then
              \state\ <= q_wait3449;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1588_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3447;
            end if;
          when q_wait3454 =>
            \$v3455\ := \$arr3399_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3451\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1588_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1578\(0 to 35) & \$1072_rest_loop668_arg\(0 to 35) & "0001" & \$v3451\;
              \state\ <= pause_setI3452;
            end if;
          when q_wait3458 =>
            \$v3459\ := \$arr3404_ptr_take\;
            if \$v3459\(0) = '1' then
              \state\ <= q_wait3458;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3456;
            end if;
          when q_wait3462 =>
            \$v3463\ := \$arr3400_ptr_take\;
            if \$v3463\(0) = '1' then
              \state\ <= q_wait3462;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= \$1603\;
              \state\ <= pause_setI3460;
            end if;
          when q_wait3470 =>
            \$v3471\ := \$arr3399_ptr_take\;
            if \$v3471\(0) = '1' then
              \state\ <= q_wait3470;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1614_t\));
              \state\ <= pause_getI3468;
            end if;
          when q_wait3476 =>
            \$v3477\ := \$arr3400_ptr_take\;
            if \$v3477\(0) = '1' then
              \state\ <= q_wait3476;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3474;
            end if;
          when q_wait3485 =>
            \$v3486\ := \$arr3399_ptr_take\;
            if \$v3486\(0) = '1' then
              \state\ <= q_wait3485;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1626_t\));
              \state\ <= pause_getI3483;
            end if;
          when q_wait3491 =>
            \$v3492\ := \$arr3400_ptr_take\;
            if \$v3492\(0) = '1' then
              \state\ <= q_wait3491;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3489;
            end if;
          when q_wait3495 =>
            \$v3496\ := \$arr3399_ptr_take\;
            if \$v3496\(0) = '1' then
              \state\ <= q_wait3495;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1635\));
              \state\ <= pause_getI3493;
            end if;
          when q_wait3499 =>
            \$v3500\ := \$arr3400_ptr_take\;
            if \$v3500\(0) = '1' then
              \state\ <= q_wait3499;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3497;
            end if;
          when q_wait3506 =>
            \$v3507\ := \$arr3399_ptr_take\;
            if \$v3507\(0) = '1' then
              \state\ <= q_wait3506;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3501\ := eclat_add(\$1072_rest_loop668_arg\(100 to 131) & "00000000000000000000000000000001");
              \$v3502\ := "00000000000000000000000000000000";
              \$v3503\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1072_rest_loop668_arg\(68 to 99)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3501\ & "0001" & \$v3502\ & "0001" & \$v3503\;
              \state\ <= pause_setI3504;
            end if;
          when q_wait3510 =>
            \$v3511\ := \$arr3400_ptr_take\;
            if \$v3511\(0) = '1' then
              \state\ <= q_wait3510;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= \$1569\;
              \state\ <= pause_setI3508;
            end if;
          when q_wait3514 =>
            \$v3515\ := \$arr3404_ptr_take\;
            if \$v3515\(0) = '1' then
              \state\ <= q_wait3514;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3512;
            end if;
          when q_wait3518 =>
            \$v3519\ := \$arr3404_ptr_take\;
            if \$v3519\(0) = '1' then
              \state\ <= q_wait3518;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1571_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3516;
            end if;
          when q_wait3522 =>
            \$v3523\ := \$arr3399_ptr_take\;
            if \$v3523\(0) = '1' then
              \state\ <= q_wait3522;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1571_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1570\;
              \state\ <= pause_setI3520;
            end if;
          when q_wait3526 =>
            \$v3527\ := \$arr3404_ptr_take\;
            if \$v3527\(0) = '1' then
              \state\ <= q_wait3526;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3524;
            end if;
          when q_wait3531 =>
            \$v3532\ := \$arr3400_ptr_take\;
            if \$v3532\(0) = '1' then
              \state\ <= q_wait3531;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3529;
            end if;
          when q_wait3536 =>
            \$v3537\ := \$arr3404_ptr_take\;
            if \$v3537\(0) = '1' then
              \state\ <= q_wait3536;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3534;
            end if;
          when q_wait3540 =>
            \$v3541\ := \$arr3404_ptr_take\;
            if \$v3541\(0) = '1' then
              \state\ <= q_wait3540;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= eclat_sub(\$1504_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3538;
            end if;
          when q_wait3545 =>
            \$v3546\ := \$arr3399_ptr_take\;
            if \$v3546\(0) = '1' then
              \state\ <= q_wait3545;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3542\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1504_i\ & "00000000000000000000000000000001")));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1494\(0 to 35) & \$1073_loop667_arg\(32 to 67) & "0001" & \$v3542\;
              \state\ <= pause_setI3543;
            end if;
          when q_wait3549 =>
            \$v3550\ := \$arr3404_ptr_take\;
            if \$v3550\(0) = '1' then
              \state\ <= q_wait3549;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr\ <= 0;
              \state\ <= pause_getI3547;
            end if;
          when q_wait3553 =>
            \$v3554\ := \$arr3400_ptr_take\;
            if \$v3554\(0) = '1' then
              \state\ <= q_wait3553;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= \$1519\;
              \state\ <= pause_setI3551;
            end if;
          when q_wait3561 =>
            \$v3562\ := \$arr3399_ptr_take\;
            if \$v3562\(0) = '1' then
              \state\ <= q_wait3561;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1530_t\));
              \state\ <= pause_getI3559;
            end if;
          when q_wait3567 =>
            \$v3568\ := \$arr3400_ptr_take\;
            if \$v3568\(0) = '1' then
              \state\ <= q_wait3567;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3565;
            end if;
          when q_wait3576 =>
            \$v3577\ := \$arr3399_ptr_take\;
            if \$v3577\(0) = '1' then
              \state\ <= q_wait3576;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1542_t\));
              \state\ <= pause_getI3574;
            end if;
          when q_wait3582 =>
            \$v3583\ := \$arr3400_ptr_take\;
            if \$v3583\(0) = '1' then
              \state\ <= q_wait3582;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3580;
            end if;
          when q_wait3586 =>
            \$v3587\ := \$arr3399_ptr_take\;
            if \$v3587\(0) = '1' then
              \state\ <= q_wait3586;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1551\));
              \state\ <= pause_getI3584;
            end if;
          when q_wait3590 =>
            \$v3591\ := \$arr3400_ptr_take\;
            if \$v3591\(0) = '1' then
              \state\ <= q_wait3590;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3588;
            end if;
          when q_wait3603 =>
            \$v3604\ := \$arr3399_ptr_take\;
            if \$v3604\(0) = '1' then
              \state\ <= q_wait3603;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
              \state\ <= pause_getI3601;
            end if;
          when q_wait3612 =>
            \$v3613\ := \$arr3400_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3610;
            end if;
          when q_wait3616 =>
            \$v3617\ := \$arr3400_ptr_take\;
            if \$v3617\(0) = '1' then
              \state\ <= q_wait3616;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= \$1395\;
              \state\ <= pause_setI3614;
            end if;
          when q_wait3623 =>
            \$v3624\ := \$arr3401_ptr_take\;
            if \$v3624\(0) = '1' then
              \state\ <= q_wait3623;
            else
              \$arr3401_ptr_take\(0) := '1';
              \$arr3401_ptr_write\ <= 0;
              \$arr3401_write_request\ <= '1';
              \$arr3401_write\ <= \$1404\;
              \state\ <= pause_setI3621;
            end if;
          when q_wait3631 =>
            \$v3632\ := \$arr3399_ptr_take\;
            if \$v3632\(0) = '1' then
              \state\ <= q_wait3631;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1414_t\));
              \state\ <= pause_getI3629;
            end if;
          when q_wait3639 =>
            \$v3640\ := \$arr3399_ptr_take\;
            if \$v3640\(0) = '1' then
              \state\ <= q_wait3639;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
              \state\ <= pause_getI3637;
            end if;
          when q_wait3648 =>
            \$v3649\ := \$arr3399_ptr_take\;
            if \$v3649\(0) = '1' then
              \state\ <= q_wait3648;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1429_t\));
              \state\ <= pause_getI3646;
            end if;
          when q_wait3654 =>
            \$v3655\ := \$arr3399_ptr_take\;
            if \$v3655\(0) = '1' then
              \state\ <= q_wait3654;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1490\;
              \state\ <= pause_setI3652;
            end if;
          when q_wait3658 =>
            \$v3659\ := \$arr3400_ptr_take\;
            if \$v3659\(0) = '1' then
              \state\ <= q_wait3658;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3656;
            end if;
          when q_wait3662 =>
            \$v3663\ := \$arr3399_ptr_take\;
            if \$v3663\(0) = '1' then
              \state\ <= q_wait3662;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \state\ <= pause_getI3660;
            end if;
          when q_wait3666 =>
            \$v3667\ := \$arr3399_ptr_take\;
            if \$v3667\(0) = '1' then
              \state\ <= q_wait3666;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1443\;
              \state\ <= pause_setI3664;
            end if;
          when q_wait3671 =>
            \$v3672\ := \$arr3399_ptr_take\;
            if \$v3672\(0) = '1' then
              \state\ <= q_wait3671;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1446_t\));
              \state\ <= pause_getI3669;
            end if;
          when q_wait3678 =>
            \$v3679\ := \$arr3399_ptr_take\;
            if \$v3679\(0) = '1' then
              \state\ <= q_wait3678;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1454_t\));
              \state\ <= pause_getI3676;
            end if;
          when q_wait3684 =>
            \$v3685\ := \$arr3399_ptr_take\;
            if \$v3685\(0) = '1' then
              \state\ <= q_wait3684;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1073_loop667_arg\(140 to 171)));
              \state\ <= pause_getI3682;
            end if;
          when q_wait3698 =>
            \$v3699\ := \$arr3399_ptr_take\;
            if \$v3699\(0) = '1' then
              \state\ <= q_wait3698;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
              \state\ <= pause_getI3696;
            end if;
          when q_wait3708 =>
            \$v3709\ := \$arr3399_ptr_take\;
            if \$v3709\(0) = '1' then
              \state\ <= q_wait3708;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1009_t\));
              \state\ <= pause_getI3706;
            end if;
          when q_wait3723 =>
            \$v3724\ := \$arr3399_ptr_take\;
            if \$v3724\(0) = '1' then
              \state\ <= q_wait3723;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1049_i\));
              \state\ <= pause_getI3721;
            end if;
          when q_wait3735 =>
            \$v3736\ := \$arr3399_ptr_take\;
            if \$v3736\(0) = '1' then
              \state\ <= q_wait3735;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1477_t\));
              \state\ <= pause_getI3733;
            end if;
          when q_wait3741 =>
            \$v3742\ := \$arr3400_ptr_take\;
            if \$v3742\(0) = '1' then
              \state\ <= q_wait3741;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3739;
            end if;
          when q_wait3750 =>
            \$v3751\ := \$arr3402_ptr_take\;
            if \$v3751\(0) = '1' then
              \state\ <= q_wait3750;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= \$1107\;
              \state\ <= pause_setI3748;
            end if;
          when q_wait3758 =>
            \$v3759\ := \$arr3399_ptr_take\;
            if \$v3759\(0) = '1' then
              \state\ <= q_wait3758;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1118_t\));
              \state\ <= pause_getI3756;
            end if;
          when q_wait3764 =>
            \$v3765\ := \$arr3402_ptr_take\;
            if \$v3765\(0) = '1' then
              \state\ <= q_wait3764;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3762;
            end if;
          when q_wait3769 =>
            \$v3770\ := \$arr3399_ptr_take\;
            if \$v3770\(0) = '1' then
              \state\ <= q_wait3769;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3766\ := "00000000000000000000000000000010";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1127\));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3766\ & \$1102\(36 to 71) & \$1102\(72 to 107);
              \state\ <= pause_setI3767;
            end if;
          when q_wait3776 =>
            \$v3777\ := \$arr3399_ptr_take\;
            if \$v3777\(0) = '1' then
              \state\ <= q_wait3776;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1138\));
              \state\ <= pause_getI3774;
            end if;
          when q_wait3784 =>
            \$v3785\ := \$arr3399_ptr_take\;
            if \$v3785\(0) = '1' then
              \state\ <= q_wait3784;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1148_t\));
              \state\ <= pause_getI3782;
            end if;
          when q_wait3790 =>
            \$v3791\ := \$arr3402_ptr_take\;
            if \$v3791\(0) = '1' then
              \state\ <= q_wait3790;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3788;
            end if;
          when q_wait3794 =>
            \$v3795\ := \$arr3402_ptr_take\;
            if \$v3795\(0) = '1' then
              \state\ <= q_wait3794;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= \$1163\;
              \state\ <= pause_setI3792;
            end if;
          when q_wait3802 =>
            \$v3803\ := \$arr3399_ptr_take\;
            if \$v3803\(0) = '1' then
              \state\ <= q_wait3802;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1174_t\));
              \state\ <= pause_getI3800;
            end if;
          when q_wait3808 =>
            \$v3809\ := \$arr3402_ptr_take\;
            if \$v3809\(0) = '1' then
              \state\ <= q_wait3808;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3806;
            end if;
          when q_wait3813 =>
            \$v3814\ := \$arr3399_ptr_take\;
            if \$v3814\(0) = '1' then
              \state\ <= q_wait3813;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3810\ := "00000000000000000000000000000001";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1183\));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3810\ & \$1158\(36 to 71) & \$1158\(72 to 107);
              \state\ <= pause_setI3811;
            end if;
          when q_wait3820 =>
            \$v3821\ := \$arr3399_ptr_take\;
            if \$v3821\(0) = '1' then
              \state\ <= q_wait3820;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1194\));
              \state\ <= pause_getI3818;
            end if;
          when q_wait3828 =>
            \$v3829\ := \$arr3399_ptr_take\;
            if \$v3829\(0) = '1' then
              \state\ <= q_wait3828;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1204_t\));
              \state\ <= pause_getI3826;
            end if;
          when q_wait3834 =>
            \$v3835\ := \$arr3402_ptr_take\;
            if \$v3835\(0) = '1' then
              \state\ <= q_wait3834;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3832;
            end if;
          when q_wait3838 =>
            \$v3839\ := \$arr3402_ptr_take\;
            if \$v3839\(0) = '1' then
              \state\ <= q_wait3838;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= \$1219\;
              \state\ <= pause_setI3836;
            end if;
          when q_wait3846 =>
            \$v3847\ := \$arr3399_ptr_take\;
            if \$v3847\(0) = '1' then
              \state\ <= q_wait3846;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1230_t\));
              \state\ <= pause_getI3844;
            end if;
          when q_wait3852 =>
            \$v3853\ := \$arr3402_ptr_take\;
            if \$v3853\(0) = '1' then
              \state\ <= q_wait3852;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3850;
            end if;
          when q_wait3857 =>
            \$v3858\ := \$arr3399_ptr_take\;
            if \$v3858\(0) = '1' then
              \state\ <= q_wait3857;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3854\ := "00000000000000000000000000000011";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1239\));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3854\ & \$1214\(36 to 71) & \$1214\(72 to 107);
              \state\ <= pause_setI3855;
            end if;
          when q_wait3864 =>
            \$v3865\ := \$arr3399_ptr_take\;
            if \$v3865\(0) = '1' then
              \state\ <= q_wait3864;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1250\));
              \state\ <= pause_getI3862;
            end if;
          when q_wait3872 =>
            \$v3873\ := \$arr3399_ptr_take\;
            if \$v3873\(0) = '1' then
              \state\ <= q_wait3872;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1260_t\));
              \state\ <= pause_getI3870;
            end if;
          when q_wait3878 =>
            \$v3879\ := \$arr3402_ptr_take\;
            if \$v3879\(0) = '1' then
              \state\ <= q_wait3878;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3876;
            end if;
          when q_wait3882 =>
            \$v3883\ := \$arr3402_ptr_take\;
            if \$v3883\(0) = '1' then
              \state\ <= q_wait3882;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= \$1275\;
              \state\ <= pause_setI3880;
            end if;
          when q_wait3890 =>
            \$v3891\ := \$arr3399_ptr_take\;
            if \$v3891\(0) = '1' then
              \state\ <= q_wait3890;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1286_t\));
              \state\ <= pause_getI3888;
            end if;
          when q_wait3896 =>
            \$v3897\ := \$arr3402_ptr_take\;
            if \$v3897\(0) = '1' then
              \state\ <= q_wait3896;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3894;
            end if;
          when q_wait3901 =>
            \$v3902\ := \$arr3399_ptr_take\;
            if \$v3902\(0) = '1' then
              \state\ <= q_wait3901;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3898\ := "00000000000000000000000000000000";
              \$arr3399_ptr_write\ <= to_integer(unsigned(\$1295\));
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3898\ & \$1270\(36 to 71) & \$1270\(72 to 107);
              \state\ <= pause_setI3899;
            end if;
          when q_wait3908 =>
            \$v3909\ := \$arr3399_ptr_take\;
            if \$v3909\(0) = '1' then
              \state\ <= q_wait3908;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1306\));
              \state\ <= pause_getI3906;
            end if;
          when q_wait3916 =>
            \$v3917\ := \$arr3399_ptr_take\;
            if \$v3917\(0) = '1' then
              \state\ <= q_wait3916;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr\ <= to_integer(unsigned(\$1316_t\));
              \state\ <= pause_getI3914;
            end if;
          when q_wait3922 =>
            \$v3923\ := \$arr3402_ptr_take\;
            if \$v3923\(0) = '1' then
              \state\ <= q_wait3922;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3920;
            end if;
          when q_wait3926 =>
            \$v3927\ := \$arr3404_ptr_take\;
            if \$v3927\(0) = '1' then
              \state\ <= q_wait3926;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= \$1325\;
              \state\ <= pause_setI3924;
            end if;
          when q_wait3930 =>
            \$v3931\ := \$arr3400_ptr_take\;
            if \$v3931\(0) = '1' then
              \state\ <= q_wait3930;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr\ <= 0;
              \state\ <= pause_getI3928;
            end if;
          when q_wait3934 =>
            \$v3935\ := \$arr3401_ptr_take\;
            if \$v3935\(0) = '1' then
              \state\ <= q_wait3934;
            else
              \$arr3401_ptr_take\(0) := '1';
              \$arr3401_ptr_write\ <= 0;
              \$arr3401_write_request\ <= '1';
              \$arr3401_write\ <= \$1326\;
              \state\ <= pause_setI3932;
            end if;
          when q_wait3938 =>
            \$v3939\ := \$arr3402_ptr_take\;
            if \$v3939\(0) = '1' then
              \state\ <= q_wait3938;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3936;
            end if;
          when q_wait3942 =>
            \$v3943\ := \$arr3399_ptr_take\;
            if \$v3943\(0) = '1' then
              \state\ <= q_wait3942;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$arr3399_ptr_write\ <= 0;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= \$1327\;
              \state\ <= pause_setI3940;
            end if;
          when q_wait3948 =>
            \$v3949\ := \$arr3402_ptr_take\;
            if \$v3949\(0) = '1' then
              \state\ <= q_wait3948;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3946;
            end if;
          when q_wait3952 =>
            \$v3953\ := \$arr3404_ptr_take\;
            if \$v3953\(0) = '1' then
              \state\ <= q_wait3952;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= \$1337\;
              \state\ <= pause_setI3950;
            end if;
          when q_wait3956 =>
            \$v3957\ := \$arr3402_ptr_take\;
            if \$v3957\(0) = '1' then
              \state\ <= q_wait3956;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr\ <= 0;
              \state\ <= pause_getI3954;
            end if;
          when q_wait3960 =>
            \$v3961\ := \$arr3402_ptr_take\;
            if \$v3961\(0) = '1' then
              \state\ <= q_wait3960;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= "00000000000000000000000000000011";
              \state\ <= pause_setI3958;
            end if;
          when q_wait3967 =>
            \$v3968\ := \$arr3399_ptr_take\;
            if \$v3968\(0) = '1' then
              \state\ <= q_wait3967;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3962\ := "00000000000000000000000000000001";
              \$v3963\ := "00000000000000000000000000000010";
              \$v3964\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 3;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0010" & \$v3962\ & "0010" & \$v3963\ & "0001" & \$v3964\;
              \state\ <= pause_setI3965;
            end if;
          when q_wait3974 =>
            \$v3975\ := \$arr3399_ptr_take\;
            if \$v3975\(0) = '1' then
              \state\ <= q_wait3974;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3969\ := "00000000000000000000000000000000";
              \$v3970\ := "00000000000000000000000000000000";
              \$v3971\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 2;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3969\ & "0001" & \$v3970\ & "0001" & \$v3971\;
              \state\ <= pause_setI3972;
            end if;
          when q_wait3981 =>
            \$v3982\ := \$arr3399_ptr_take\;
            if \$v3982\(0) = '1' then
              \state\ <= q_wait3981;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3976\ := "00000000000000000000000000000000";
              \$v3977\ := "00000000000000000000000000000000";
              \$v3978\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 1;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3976\ & "0001" & \$v3977\ & "0001" & \$v3978\;
              \state\ <= pause_setI3979;
            end if;
          when q_wait3988 =>
            \$v3989\ := \$arr3399_ptr_take\;
            if \$v3989\(0) = '1' then
              \state\ <= q_wait3988;
            else
              \$arr3399_ptr_take\(0) := '1';
              \$v3983\ := "00000000000000000000000000000000";
              \$v3984\ := "00000000000000000000000000000000";
              \$v3985\ := "00000000000000000000000000000101";
              \$arr3399_ptr_write\ <= 0;
              \$arr3399_write_request\ <= '1';
              \$arr3399_write\ <= "0001" & \$v3983\ & "0001" & \$v3984\ & "0001" & \$v3985\;
              \state\ <= pause_setI3986;
            end if;
          when q_wait3992 =>
            \$v3993\ := \$arr3405_ptr_take\;
            if \$v3993\(0) = '1' then
              \state\ <= q_wait3992;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 5;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI3990;
            end if;
          when q_wait3996 =>
            \$v3997\ := \$arr3405_ptr_take\;
            if \$v3997\(0) = '1' then
              \state\ <= q_wait3996;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 4;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI3994;
            end if;
          when q_wait4000 =>
            \$v4001\ := \$arr3405_ptr_take\;
            if \$v4001\(0) = '1' then
              \state\ <= q_wait4000;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 3;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI3998;
            end if;
          when q_wait4004 =>
            \$v4005\ := \$arr3405_ptr_take\;
            if \$v4005\(0) = '1' then
              \state\ <= q_wait4004;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 2;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4002;
            end if;
          when q_wait4008 =>
            \$v4009\ := \$arr3405_ptr_take\;
            if \$v4009\(0) = '1' then
              \state\ <= q_wait4008;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 1;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI4006;
            end if;
          when q_wait4012 =>
            \$v4013\ := \$arr3405_ptr_take\;
            if \$v4013\(0) = '1' then
              \state\ <= q_wait4012;
            else
              \$arr3405_ptr_take\(0) := '1';
              \$arr3405_ptr_write\ <= 0;
              \$arr3405_write_request\ <= '1';
              \$arr3405_write\ <= X"000000" & X"14";
              \state\ <= pause_setI4010;
            end if;
          when q_wait4016 =>
            \$v4017\ := \$arr3404_ptr_take\;
            if \$v4017\(0) = '1' then
              \state\ <= q_wait4016;
            else
              \$arr3404_ptr_take\(0) := '1';
              \$arr3404_ptr_write\ <= 0;
              \$arr3404_write_request\ <= '1';
              \$arr3404_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4014;
            end if;
          when q_wait4020 =>
            \$v4021\ := \$arr3403_ptr_take\;
            if \$v4021\(0) = '1' then
              \state\ <= q_wait4020;
            else
              \$arr3403_ptr_take\(0) := '1';
              \$arr3403_ptr_write\ <= 0;
              \$arr3403_write_request\ <= '1';
              \$arr3403_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4018;
            end if;
          when q_wait4024 =>
            \$v4025\ := \$arr3402_ptr_take\;
            if \$v4025\(0) = '1' then
              \state\ <= q_wait4024;
            else
              \$arr3402_ptr_take\(0) := '1';
              \$arr3402_ptr_write\ <= 0;
              \$arr3402_write_request\ <= '1';
              \$arr3402_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4022;
            end if;
          when q_wait4028 =>
            \$v4029\ := \$arr3400_ptr_take\;
            if \$v4029\(0) = '1' then
              \state\ <= q_wait4028;
            else
              \$arr3400_ptr_take\(0) := '1';
              \$arr3400_ptr_write\ <= 0;
              \$arr3400_write_request\ <= '1';
              \$arr3400_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI4026;
            end if;
          when q_wait4032 =>
            \$v4033\ := \$arr3401_ptr_take\;
            if \$v4033\(0) = '1' then
              \state\ <= q_wait4032;
            else
              \$arr3401_ptr_take\(0) := '1';
              \$arr3401_ptr_write\ <= 0;
              \$arr3401_write_request\ <= '1';
              \$arr3401_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4030;
            end if;
          when compute3408 =>
            rdy3407 := eclat_false;
            \$v4033\ := \$arr3401_ptr_take\;
            if \$v4033\(0) = '1' then
              \state\ <= q_wait4032;
            else
              \$arr3401_ptr_take\(0) := '1';
              \$arr3401_ptr_write\ <= 0;
              \$arr3401_write_request\ <= '1';
              \$arr3401_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI4030;
            end if;
          end case;
          
          result <= result3406;
          rdy <= rdy3407;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
