-- code generated from the following source code:
--   ../RibbitVm/fail.ecl
--   ../RibbitVm/vm.ecl
--
-- with the following command:
--
--    ./eclat ../RibbitVm/fail.ecl ../RibbitVm/vm.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute3246, \$1046_list_tail618\, \$1047_get_int621\, \$1049_rest_loop649\, \$1050_loop648\, \$1085_show_rib6123223\, \$1102_forever6703195\, \$1114_forever6703224\, \$1124_forever6703225\, \$1132_forever6703226\, \$1137_print_value5913227\, \$1147_forever6703228\, \$1164_forever6703229\, \$1172_forever6703230\, \$1178_loop6503231\, \$1187_forever6703214\, \$1195_forever6703218\, \$1229_forever6703232\, \$1239_forever6703233\, \$1248_forever6703234\, \$1260_forever6703235\, \$1313_forever6703219\, \$1323_forever6703220\, \$1332_forever6703221\, \$1344_forever6703222\, \$1383_forever6703196\, \$1398_forever6703197\, \$369_forever6703193\, \$369_forever6703194\, \$369_forever6703195\, \$369_forever6703216\, \$409_show_rib6123215\, \$409_show_rib6123217\, pause_getI3251, pause_getI3259, pause_getI3269, pause_getI3273, pause_getI3277, pause_getI3281, pause_getI3294, pause_getI3306, pause_getI3312, pause_getI3321, pause_getI3327, pause_getI3331, pause_getI3335, pause_getI3350, pause_getI3362, pause_getI3367, pause_getI3372, pause_getI3385, pause_getI3397, pause_getI3403, pause_getI3412, pause_getI3418, pause_getI3422, pause_getI3426, pause_getI3439, pause_getI3448, pause_getI3467, pause_getI3475, pause_getI3484, pause_getI3494, pause_getI3498, pause_getI3507, pause_getI3514, pause_getI3520, pause_getI3534, pause_getI3544, pause_getI3559, pause_getI3571, pause_getI3577, pause_getII3252, pause_getII3260, pause_getII3270, pause_getII3274, pause_getII3278, pause_getII3282, pause_getII3295, pause_getII3307, pause_getII3313, pause_getII3322, pause_getII3328, pause_getII3332, pause_getII3336, pause_getII3351, pause_getII3363, pause_getII3368, pause_getII3373, pause_getII3386, pause_getII3398, pause_getII3404, pause_getII3413, pause_getII3419, pause_getII3423, pause_getII3427, pause_getII3440, pause_getII3449, pause_getII3468, pause_getII3476, pause_getII3485, pause_getII3495, pause_getII3499, pause_getII3508, pause_getII3515, pause_getII3521, pause_getII3535, pause_getII3545, pause_getII3560, pause_getII3572, pause_getII3578, pause_setI3265, pause_setI3285, pause_setI3290, pause_setI3298, pause_setI3342, pause_setI3346, pause_setI3354, pause_setI3358, pause_setI3376, pause_setI3381, pause_setI3389, pause_setI3452, pause_setI3459, pause_setI3490, pause_setI3502, pause_setI3586, pause_setI3590, pause_setI3594, pause_setI3598, pause_setI3602, pause_setI3606, pause_setI3610, pause_setI3614, pause_setI3618, pause_setI3622, pause_setI3626, pause_setII3266, pause_setII3286, pause_setII3291, pause_setII3299, pause_setII3343, pause_setII3347, pause_setII3355, pause_setII3359, pause_setII3377, pause_setII3382, pause_setII3390, pause_setII3453, pause_setII3460, pause_setII3491, pause_setII3503, pause_setII3587, pause_setII3591, pause_setII3595, pause_setII3599, pause_setII3603, pause_setII3607, pause_setII3611, pause_setII3615, pause_setII3619, pause_setII3623, pause_setII3627, q_wait3253, q_wait3261, q_wait3267, q_wait3271, q_wait3275, q_wait3279, q_wait3283, q_wait3287, q_wait3292, q_wait3296, q_wait3300, q_wait3308, q_wait3314, q_wait3323, q_wait3329, q_wait3333, q_wait3337, q_wait3344, q_wait3348, q_wait3352, q_wait3356, q_wait3360, q_wait3364, q_wait3369, q_wait3374, q_wait3378, q_wait3383, q_wait3387, q_wait3391, q_wait3399, q_wait3405, q_wait3414, q_wait3420, q_wait3424, q_wait3428, q_wait3441, q_wait3450, q_wait3454, q_wait3461, q_wait3469, q_wait3477, q_wait3486, q_wait3492, q_wait3496, q_wait3500, q_wait3504, q_wait3509, q_wait3516, q_wait3522, q_wait3536, q_wait3546, q_wait3561, q_wait3573, q_wait3579, q_wait3588, q_wait3592, q_wait3596, q_wait3600, q_wait3604, q_wait3608, q_wait3612, q_wait3616, q_wait3620, q_wait3624, q_wait3628);
  signal \state\: t_state;
  type array_value_32 is array (natural range <>) of value(0 to 31);
  type array_value_108 is array (natural range <>) of value(0 to 107);
  signal arr3236 : array_value_32(0 to 8999) := (others => (others => '0'));
  signal \$arr3236_value\ : value(0 to 31);
  signal \$arr3236_ptr\ : natural range 0 to 8999;
  signal \$arr3236_ptr_write\ : natural range 0 to 8999;
  signal \$arr3236_write\ : value(0 to 31);
  signal \$arr3236_write_request\ : std_logic := '0';
  signal arr3237 : array_value_108(0 to 8999) := (others => (others => '0'));
  signal \$arr3237_value\ : value(0 to 107);
  signal \$arr3237_ptr\ : natural range 0 to 8999;
  signal \$arr3237_ptr_write\ : natural range 0 to 8999;
  signal \$arr3237_write\ : value(0 to 107);
  signal \$arr3237_write_request\ : std_logic := '0';
  signal arr3238 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3238_value\ : value(0 to 31);
  signal \$arr3238_ptr\ : natural range 0 to 0;
  signal \$arr3238_ptr_write\ : natural range 0 to 0;
  signal \$arr3238_write\ : value(0 to 31);
  signal \$arr3238_write_request\ : std_logic := '0';
  signal arr3239 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3239_value\ : value(0 to 31);
  signal \$arr3239_ptr\ : natural range 0 to 0;
  signal \$arr3239_ptr_write\ : natural range 0 to 0;
  signal \$arr3239_write\ : value(0 to 31);
  signal \$arr3239_write_request\ : std_logic := '0';
  signal arr3240 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3240_value\ : value(0 to 31);
  signal \$arr3240_ptr\ : natural range 0 to 0;
  signal \$arr3240_ptr_write\ : natural range 0 to 0;
  signal \$arr3240_write\ : value(0 to 31);
  signal \$arr3240_write_request\ : std_logic := '0';
  signal arr3241 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3241_value\ : value(0 to 31);
  signal \$arr3241_ptr\ : natural range 0 to 0;
  signal \$arr3241_ptr_write\ : natural range 0 to 0;
  signal \$arr3241_write\ : value(0 to 31);
  signal \$arr3241_write_request\ : std_logic := '0';
  signal arr3242 : array_value_32(0 to 0) := (others => (others => '0'));
  signal \$arr3242_value\ : value(0 to 31);
  signal \$arr3242_ptr\ : natural range 0 to 0;
  signal \$arr3242_ptr_write\ : natural range 0 to 0;
  signal \$arr3242_write\ : value(0 to 31);
  signal \$arr3242_write_request\ : std_logic := '0';
  signal arr3243 : array_value_32(0 to 5) := (others => (others => '0'));
  signal \$arr3243_value\ : value(0 to 31);
  signal \$arr3243_ptr\ : natural range 0 to 5;
  signal \$arr3243_ptr_write\ : natural range 0 to 5;
  signal \$arr3243_write\ : value(0 to 31);
  signal \$arr3243_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3236_write_request\ = '1' then
                    arr3236(\$arr3236_ptr_write\) <= \$arr3236_write\;
                  else
                   \$arr3236_value\ <= arr3236(\$arr3236_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3237_write_request\ = '1' then
                    arr3237(\$arr3237_ptr_write\) <= \$arr3237_write\;
                  else
                   \$arr3237_value\ <= arr3237(\$arr3237_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3238_write_request\ = '1' then
                    arr3238(\$arr3238_ptr_write\) <= \$arr3238_write\;
                  else
                   \$arr3238_value\ <= arr3238(\$arr3238_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3239_write_request\ = '1' then
                    arr3239(\$arr3239_ptr_write\) <= \$arr3239_write\;
                  else
                   \$arr3239_value\ <= arr3239(\$arr3239_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3240_write_request\ = '1' then
                    arr3240(\$arr3240_ptr_write\) <= \$arr3240_write\;
                  else
                   \$arr3240_value\ <= arr3240(\$arr3240_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3241_write_request\ = '1' then
                    arr3241(\$arr3241_ptr_write\) <= \$arr3241_write\;
                  else
                   \$arr3241_value\ <= arr3241(\$arr3241_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3242_write_request\ = '1' then
                    arr3242(\$arr3242_ptr_write\) <= \$arr3242_write\;
                  else
                   \$arr3242_value\ <= arr3242(\$arr3242_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr3243_write_request\ = '1' then
                    arr3243(\$arr3243_ptr_write\) <= \$arr3243_write\;
                  else
                   \$arr3243_value\ <= arr3243(\$arr3243_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$v3583\, \$v3435\, \$v3325\, \$v3257\, 
               \$1137_print_value5913227_arg\, \$v3548\, \$1299\, \$v3530\, 
               \$1177\, \$v3479\, \$v3526\, \$v3575\, \$v3416\, \$1234\, 
               \$1318\, \$v3394\, \$1107\, \$v3471\, \$v3568\, \$v3249\, 
               \$v3457\, \$1289\, \$v3303\, \$v3540\, \$v3565\, 
               \$1178_loop6503231_arg\, \$1158\, \$1402\, \$v3310\, \$v3318\, 
               \$v3445\, \$v3511\, \$1255\, \$v3464\, \$v3563\, \$1339\, 
               \$v3518\, \$v3431\, \$1243\, \$v3443\, \$1136\, \$v3401\, 
               \$v3481\, \$1215\, \$1181_tag\, \$1253\, 
               \$1178_loop6503231_result\, \$1119\, \$v3538\, \$v3551\, 
               \$1152_k\, \$1327\, \$v3409\, \$1159\, \$1337\, \$1205\, 
               \$v3555\, \$v405\, \$v3488\ : value(0 to 35) := (others => '0');
      variable \$1391\, \$1364\, \$1046_list_tail618_arg\, \$1370\ : value(0 to 63) := (others => '0');
      variable \$1049_rest_loop649_arg\ : value(0 to 131) := (others => '0');
      variable \$v3480\, \$v3432\, \$v3569\, \$v3250\, \$v3566\, \$v3489\, 
               \$v3539\, \$v3417\, \$v3304\, \$v3576\, \$v3552\, \$v3311\, 
               \$v3564\, \$v3549\, \$v3519\, \$v3482\, \$v3326\, \$v3584\, 
               \$v3258\, \$v3402\, \$v3436\, \$v3458\, \$v3444\, \$v3512\, 
               \$v3472\, \$v3319\, \$v3527\, \$v3556\, \$v3410\, \$v3541\, 
               \$v3465\, \$v3446\, \$v3531\, \$v3395\ : value(0 to 3) := (others => '0');
      variable \$1137_print_value5913227_result\, \$v3371\, 
               \$409_show_rib6123215_result\, \$v3567\, \$v3609\, \$v3574\, 
               result3244, \$v3375\, \$1151\, \$v3297\, \$v3268\, \$1309\, 
               \$v3589\, \$v3580\, \$v3334\, \$v3447\, \$v3349\, \$v3254\, 
               \$v3593\, \$v3553\, \$881\, \$v3264\, rdy3245, \$v3497\, 
               \$409_show_rib6123217_result\, \$v3621\, \$v3301\, \$v3262\, 
               \$1096\, \$v3415\, \$v3505\, \$v3597\, \$v3617\, \$v3288\, 
               \$v3542\, \$v3406\, \$v3407\, \$v3510\, \$v3421\, \$v3293\, 
               \$v3315\, \$v3384\, \$v3442\, \$v3316\, \$v3462\, 
               \$1085_show_rib6123223_result\, \$v3309\, \$1379\, \$v3338\, 
               \$v3276\, \$v3284\, \$v3400\, \$v3517\, \$v3433\, \$v3537\, 
               \$v3629\, \$v3263\, \$v3501\, \$v3255\, \$1225\, \$v3605\, 
               \$v3353\, \$v3429\, \$v3379\, \$v3528\, \$v3493\, \$v3370\, 
               \$v3280\, \$v3523\, \$v3601\, \$v3365\, \$v3357\, \$v3324\, 
               \$v3345\, \$v3361\, \$v3392\, \$v3625\, \$v3470\, \$v3425\, 
               \$v3455\, \$v3562\, \$v3451\, \$v3330\, \$v3585\, \$v3581\, 
               \$v3547\, \$v3272\, \$v3388\, \$v3478\, \$v3487\, \$v3613\ : value(0 to 0) := (others => '0');
      variable \$1050_loop648_arg\ : value(0 to 171) := (others => '0');
      variable \$1157\, \$v2774\, \$1404\, \$1208\, \$1292\, \$v2783\, 
               \$1153\, \$v2778\, \$1387\, \$v2808\, \$v3173\, \$v3160\, 
               \$1200\, \$v2834\, \$v2787\, \$v2804\, \$1284\, \$v2847\, 
               \$v2843\, \$v2830\, \$1204\ : value(0 to 107) := (others => '0');
      variable \$409_show_rib6123217_arg\, \$1084\, 
               \$409_show_rib6123215_arg\, \$1085_show_rib6123223_arg\ : value(0 to 99) := (others => '0');
      variable \$v3411\, \$v3570\, \$1191_t\, \$879_i\, \$1128_t\, \$1217\, 
               \$v3532\, \$1097\, \$1371\, \$v3533\, \$v3554\, \$1030_i\, 
               \$1291\, \$v3408\, \$1328_t\, \$1352_x\, \$v3463\, \$977_t\, 
               \$v3513\, \$1120_i\, \$1265\, \$v3430\, \$v3506\, \$v3305\, 
               \$1168_t\, \$1285_i\, \$882\, \$v3550\, \$1372\, \$1365\, 
               \$v3437\, \$v3456\, \$v3473\, \$v3289\, \$v3320\, \$v3466\, 
               \$1256_t\, \$v3524\, \$v3339\, \$v3317\, \$1244_t\, \$1108\, 
               \$1348\, \$v3340\, \$1199\, \$1362_x\, \$1302_i\, \$v3302\, 
               \$1317\, \$1094_i\, \$1109\, \$1218_i\, \$1252\, \$1143_t\, 
               \$v3341\, \$1026_i\, \$v3483\, \$v3434\, \$1367_c\, \$1349\, 
               \$v3396\, \$1283\, \$v3558\, \$1140_t\, \$1336\, \$1110_i\, 
               \$1369\, \$v3380\, \$v3247\, \$1319_i\, \$1301\, \$1264\, 
               \$1047_get_int621_arg\, \$1118\, \$1392\, \$v3557\, \$v3525\, 
               \$v3529\, \$1142_i\, \$1160_t\, \$v3474\, \$v3256\, \$1394_i\, 
               \$1340_t\, \$v3393\, \$v3366\, \$1098_i\, \$1233\, \$v3543\, 
               \$v3582\, \$1235_i\, \$1206\, \$v3438\, \$v3248\ : value(0 to 31) := (others => '0');
      variable \$1298\, \$1214\ : value(0 to 67) := (others => '0');
      variable \$arr3236_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3237_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3238_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3239_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3240_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3241_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3242_ptr_take\ : value(0 to 0) := "0";
      variable \$arr3243_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v3488\); default_zero(\$v405\); 
          default_zero(\$v3555\); default_zero(\$v3613\); 
          default_zero(\$v3395\); default_zero(\$1370\); 
          default_zero(\$v3248\); default_zero(\$v3438\); 
          default_zero(\$1206\); default_zero(\$1235_i\); 
          default_zero(\$1205\); default_zero(\$v3582\); 
          default_zero(\$v3487\); default_zero(\$v3543\); 
          default_zero(\$1337\); default_zero(\$v3478\); 
          default_zero(\$1085_show_rib6123223_arg\); default_zero(\$1233\); 
          default_zero(\$1098_i\); default_zero(\$v3388\); 
          default_zero(\$1204\); default_zero(\$v3366\); 
          default_zero(\$v3272\); default_zero(\$v3393\); 
          default_zero(\$1340_t\); default_zero(\$1394_i\); 
          default_zero(\$v3547\); default_zero(\$v3581\); 
          default_zero(\$v3585\); default_zero(\$v3256\); 
          default_zero(\$v3330\); default_zero(\$v3531\); 
          default_zero(\$v2830\); default_zero(\$v3474\); 
          default_zero(\$v3451\); default_zero(\$1159\); 
          default_zero(\$v3562\); default_zero(\$v2843\); 
          default_zero(\$1160_t\); default_zero(\$1142_i\); 
          default_zero(\$v3455\); default_zero(\$v3409\); 
          default_zero(\$v3446\); default_zero(\$v3425\); 
          default_zero(\$v3529\); default_zero(\$409_show_rib6123215_arg\); 
          default_zero(\$v2847\); default_zero(\$v3470\); 
          default_zero(\$v3465\); default_zero(\$v3625\); 
          default_zero(\$1327\); default_zero(\$v3392\); 
          default_zero(\$v3361\); default_zero(\$v3345\); 
          default_zero(\$v3324\); default_zero(\$v3525\); 
          default_zero(\$1152_k\); default_zero(\$v3541\); 
          default_zero(\$v3410\); default_zero(\$v3551\); 
          default_zero(\$v3556\); default_zero(\$v3538\); 
          default_zero(\$v3527\); default_zero(\$v3319\); 
          default_zero(\$1084\); default_zero(\$1284\); 
          default_zero(\$v3472\); default_zero(\$1119\); 
          default_zero(\$v3557\); default_zero(\$1392\); 
          default_zero(\$1178_loop6503231_result\); default_zero(\$v3357\); 
          default_zero(\$1118\); default_zero(\$1047_get_int621_arg\); 
          default_zero(\$v3512\); default_zero(\$1253\); 
          default_zero(\$v3365\); default_zero(\$1264\); 
          default_zero(\$v3601\); default_zero(\$1301\); 
          default_zero(\$1319_i\); default_zero(\$1181_tag\); 
          default_zero(\$v3523\); default_zero(\$1215\); 
          default_zero(\$v3280\); default_zero(\$v3370\); 
          default_zero(\$v3493\); default_zero(\$v3528\); 
          default_zero(\$v3481\); default_zero(\$v3247\); 
          default_zero(\$v3379\); default_zero(\$v3429\); 
          default_zero(\$v3353\); default_zero(\$v3380\); 
          default_zero(\$1369\); default_zero(\$1110_i\); 
          default_zero(\$v3605\); default_zero(\$v3401\); 
          default_zero(\$1336\); default_zero(\$1136\); 
          default_zero(\$v3443\); default_zero(\$1243\); 
          default_zero(\$1140_t\); default_zero(\$1225\); 
          default_zero(\$v3255\); default_zero(\$v3558\); 
          default_zero(\$v3431\); default_zero(\$v3518\); 
          default_zero(\$1283\); default_zero(\$v3396\); 
          default_zero(\$1349\); default_zero(\$v3501\); 
          default_zero(\$v3263\); default_zero(\$1339\); 
          default_zero(\$1367_c\); default_zero(\$v3444\); 
          default_zero(\$v2804\); default_zero(\$v3434\); 
          default_zero(\$v2787\); default_zero(\$v3563\); 
          default_zero(\$v3629\); default_zero(\$v3483\); 
          default_zero(\$v3537\); default_zero(\$v3458\); 
          default_zero(\$v3464\); default_zero(\$1026_i\); 
          default_zero(\$v3436\); default_zero(\$v3341\); 
          default_zero(\$1143_t\); default_zero(\$v3402\); 
          default_zero(\$v3433\); default_zero(\$v3517\); 
          default_zero(\$v3400\); default_zero(\$v3284\); 
          default_zero(\$1050_loop648_arg\); default_zero(\$1252\); 
          default_zero(\$v3276\); default_zero(\$1218_i\); 
          default_zero(\$v3258\); default_zero(\$1109\); 
          default_zero(\$1255\); default_zero(\$1214\); 
          default_zero(\$v3338\); default_zero(\$1094_i\); 
          default_zero(\$1317\); default_zero(\$v3584\); 
          default_zero(\$v3511\); default_zero(\$1379\); 
          default_zero(\$v3445\); default_zero(\$v3326\); 
          default_zero(\$v3318\); default_zero(\$v3309\); 
          default_zero(\$1085_show_rib6123223_result\); 
          default_zero(\$v3310\); default_zero(\$v3302\); 
          default_zero(\$1402\); default_zero(\$1302_i\); 
          default_zero(\$v2834\); default_zero(\$1362_x\); 
          default_zero(\$1158\); default_zero(\$v3462\); 
          default_zero(\$v3316\); default_zero(\$v3482\); 
          default_zero(\$v3442\); default_zero(\$1200\); 
          default_zero(\$v3384\); default_zero(\$v3315\); 
          default_zero(\$v3519\); default_zero(\$1199\); 
          default_zero(\$v3160\); default_zero(\$1178_loop6503231_arg\); 
          default_zero(\$v3173\); default_zero(\$v3549\); 
          default_zero(\$v3340\); default_zero(\$v2808\); 
          default_zero(\$v3565\); default_zero(\$1348\); 
          default_zero(\$1108\); default_zero(\$v3293\); 
          default_zero(\$1244_t\); default_zero(\$v3421\); 
          default_zero(\$v3317\); default_zero(\$v3339\); 
          default_zero(\$v3524\); default_zero(\$1046_list_tail618_arg\); 
          default_zero(\$v3510\); default_zero(\$1256_t\); 
          default_zero(\$v3466\); default_zero(\$v3407\); 
          default_zero(\$v3320\); default_zero(\$v3289\); 
          default_zero(\$v3473\); default_zero(\$v3406\); 
          default_zero(\$1049_rest_loop649_arg\); default_zero(\$v3542\); 
          default_zero(\$v3456\); default_zero(\$v3437\); 
          default_zero(\$v3288\); default_zero(\$1298\); 
          default_zero(\$v3617\); default_zero(\$1365\); 
          default_zero(\$v3597\); default_zero(\$v3505\); 
          default_zero(\$v3415\); default_zero(\$1372\); 
          default_zero(\$v3540\); default_zero(\$1387\); 
          default_zero(\$v3550\); default_zero(\$1096\); 
          default_zero(\$v3262\); default_zero(\$882\); 
          default_zero(\$1285_i\); default_zero(\$v3303\); 
          default_zero(\$1168_t\); default_zero(\$1289\); 
          default_zero(\$v3305\); default_zero(\$v3301\); 
          default_zero(\$v3457\); default_zero(\$v3621\); 
          default_zero(\$409_show_rib6123217_result\); 
          default_zero(\$v3249\); default_zero(\$v3568\); 
          default_zero(\$v3471\); default_zero(\$v3564\); 
          default_zero(\$v3506\); default_zero(\$v3497\); 
          default_zero(rdy3245); default_zero(\$v3264\); 
          default_zero(\$v3430\); default_zero(\$881\); 
          default_zero(\$1364\); default_zero(\$1391\); 
          default_zero(\$v3553\); default_zero(\$1107\); 
          default_zero(\$v3593\); default_zero(\$v3394\); 
          default_zero(\$1265\); default_zero(\$v3254\); 
          default_zero(\$1318\); default_zero(\$v3311\); 
          default_zero(\$1120_i\); default_zero(\$v3349\); 
          default_zero(\$v3552\); default_zero(\$v2778\); 
          default_zero(\$v3447\); default_zero(\$1234\); 
          default_zero(\$v3576\); default_zero(\$v3513\); 
          default_zero(\$977_t\); default_zero(\$v3334\); 
          default_zero(\$409_show_rib6123217_arg\); default_zero(\$v3463\); 
          default_zero(\$v3580\); default_zero(\$1352_x\); 
          default_zero(\$v3416\); default_zero(\$v3575\); 
          default_zero(\$v3589\); default_zero(\$1309\); 
          default_zero(\$1328_t\); default_zero(\$v3408\); 
          default_zero(\$v3526\); default_zero(\$v3479\); 
          default_zero(\$1177\); default_zero(\$1153\); 
          default_zero(\$v3268\); default_zero(\$v3297\); 
          default_zero(\$1291\); default_zero(\$v3530\); 
          default_zero(\$1151\); default_zero(\$1299\); 
          default_zero(\$v3304\); default_zero(\$v3375\); 
          default_zero(\$1030_i\); default_zero(result3244); 
          default_zero(\$v3554\); default_zero(\$v3574\); 
          default_zero(\$v3609\); default_zero(\$v3533\); 
          default_zero(\$v2783\); default_zero(\$1292\); 
          default_zero(\$v3567\); 
          default_zero(\$409_show_rib6123215_result\); 
          default_zero(\$v3548\); default_zero(\$v3371\); 
          default_zero(\$1371\); default_zero(\$1208\); 
          default_zero(\$1404\); default_zero(\$v3417\); 
          default_zero(\$1097\); default_zero(\$v2774\); 
          default_zero(\$v3539\); default_zero(\$v3532\); 
          default_zero(\$1157\); default_zero(\$v3489\); 
          default_zero(\$1217\); default_zero(\$v3566\); 
          default_zero(\$1128_t\); 
          default_zero(\$1137_print_value5913227_result\); 
          default_zero(\$1137_print_value5913227_arg\); 
          default_zero(\$879_i\); default_zero(\$1191_t\); 
          default_zero(\$v3257\); default_zero(\$v3570\); 
          default_zero(\$v3325\); default_zero(\$v3250\); 
          default_zero(\$v3569\); default_zero(\$v3435\); 
          default_zero(\$v3432\); default_zero(\$v3583\); 
          default_zero(\$v3480\); default_zero(\$v3411\); 
          rdy <= "1";
          rdy3245 := "0";
          \state\ <= compute3246;
          
        else if run = '1' then
          case \state\ is
          when \$1046_list_tail618\ =>
            \$v3263\ := eclat_eq("00000000000000000000000000000000" & \$1046_list_tail618_arg\(32 to 63));
            if \$v3263\(0) = '1' then
              \$v3247\ := \$1046_list_tail618_arg\(0 to 31);
              
              \state\ <= \$1046_list_tail618\;
            else
              \$v3262\ := \$arr3237_ptr_take\;
              if \$v3262\(0) = '1' then
                \state\ <= q_wait3261;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1046_list_tail618_arg\(0 to 31)));
                \state\ <= pause_getI3259;
              end if;
            end if;
          when \$1047_get_int621\ =>
            \$v3280\ := \$arr3241_ptr_take\;
            if \$v3280\(0) = '1' then
              \state\ <= q_wait3279;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr\ <= 0;
              \state\ <= pause_getI3277;
            end if;
          when \$1049_rest_loop649\ =>
            \$v3371\ := eclat_lt("00000000000000000000000000000000" & \$1049_rest_loop649_arg\(36 to 67));
            if \$v3371\(0) = '1' then
              \$v3338\ := \$arr3238_ptr_take\;
              if \$v3338\(0) = '1' then
                \state\ <= q_wait3337;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr\ <= 0;
                \state\ <= pause_getI3335;
              end if;
            else
              \$v3370\ := \$arr3238_ptr_take\;
              if \$v3370\(0) = '1' then
                \state\ <= q_wait3369;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr\ <= 0;
                \state\ <= pause_getI3367;
              end if;
            end if;
          when \$1050_loop648\ =>
            \$v3585\ := eclat_lt("00000000000000000000000000000000" & \$1050_loop648_arg\(0 to 31));
            if \$v3585\(0) = '1' then
              \$v3429\ := \$arr3238_ptr_take\;
              if \$v3429\(0) = '1' then
                \state\ <= q_wait3428;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr\ <= 0;
                \state\ <= pause_getI3426;
              end if;
            else
              \$v3583\ := \$1050_loop648_arg\(68 to 103);
              \$v3584\ := \$v3583\(0 to 3);
              \$v3582\ := \$v3583\(4 to 35);
              case \$v3584\ is
              when "0010" =>
                \$1151\ := eclat_true;
                \$v3581\ := \$1151\;
                if \$v3581\(0) = '1' then
                  \$v3501\ := \$arr3237_ptr_take\;
                  if \$v3501\(0) = '1' then
                    \state\ <= q_wait3500;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                    \state\ <= pause_getI3498;
                  end if;
                else
                  \$v3580\ := \$arr3238_ptr_take\;
                  if \$v3580\(0) = '1' then
                    \state\ <= q_wait3579;
                  else
                    \$arr3238_ptr_take\(0) := '1';
                    \$arr3238_ptr\ <= 0;
                    \state\ <= pause_getI3577;
                  end if;
                end if;
              when others =>
                \$1151\ := eclat_false;
                \$v3581\ := \$1151\;
                if \$v3581\(0) = '1' then
                  \$v3501\ := \$arr3237_ptr_take\;
                  if \$v3501\(0) = '1' then
                    \state\ <= q_wait3500;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                    \state\ <= pause_getI3498;
                  end if;
                else
                  \$v3580\ := \$arr3238_ptr_take\;
                  if \$v3580\(0) = '1' then
                    \state\ <= q_wait3579;
                  else
                    \$arr3238_ptr_take\(0) := '1';
                    \$arr3238_ptr\ <= 0;
                    \state\ <= pause_getI3577;
                  end if;
                end if;
              end case;
            end if;
          when \$1085_show_rib6123223\ =>
            \$v3447\ := eclat_gt(\$1085_show_rib6123223_arg\(68 to 99) & \$1085_show_rib6123223_arg\(36 to 67));
            if \$v3447\(0) = '1' then
              \$v3435\ := \$1085_show_rib6123223_arg\(0 to 35);
              \$v3436\ := \$v3435\(0 to 3);
              \$v3434\ := \$v3435\(4 to 35);
              case \$v3436\ is
              when "0010" =>
                \$1096\ := eclat_true;
                \$v3433\ := \$1096\;
                if \$v3433\(0) = '1' then
                  \$1085_show_rib6123223_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \state\ <= \$1050_loop648\;
                else
                  \$v3431\ := \$1085_show_rib6123223_arg\(0 to 35);
                  \$v3432\ := \$v3431\(0 to 3);
                  \$v3430\ := \$v3431\(4 to 35);
                  case \$v3432\ is
                  when "0001" =>
                    \$1098_i\ := \$v3430\(0 to 31);
                    \$1097\ := \$1098_i\;
                    \$1085_show_rib6123223_result\ := eclat_unit;
                    eclat_print_int(\$1097\);
                    
                    \state\ <= \$1050_loop648\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$1102_forever6703195\;
                  end case;
                end if;
              when others =>
                \$1096\ := eclat_false;
                \$v3433\ := \$1096\;
                if \$v3433\(0) = '1' then
                  \$1085_show_rib6123223_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \state\ <= \$1050_loop648\;
                else
                  \$v3431\ := \$1085_show_rib6123223_arg\(0 to 35);
                  \$v3432\ := \$v3431\(0 to 3);
                  \$v3430\ := \$v3431\(4 to 35);
                  case \$v3432\ is
                  when "0001" =>
                    \$1098_i\ := \$v3430\(0 to 31);
                    \$1097\ := \$1098_i\;
                    \$1085_show_rib6123223_result\ := eclat_unit;
                    eclat_print_int(\$1097\);
                    
                    \state\ <= \$1050_loop648\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$1102_forever6703195\;
                  end case;
                end if;
              end case;
            else
              \$v3445\ := \$1085_show_rib6123223_arg\(0 to 35);
              \$v3446\ := \$v3445\(0 to 3);
              \$v3437\ := \$v3445\(4 to 35);
              case \$v3446\ is
              when "0000" =>
                \$1085_show_rib6123223_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \state\ <= \$1050_loop648\;
              when "0001" =>
                \$1094_i\ := \$v3437\(0 to 31);
                \$1085_show_rib6123223_result\ := eclat_unit;
                eclat_print_int(\$1094_i\);
                
                \state\ <= \$1050_loop648\;
              when "0010" =>
                \$v3443\ := \$1085_show_rib6123223_arg\(0 to 35);
                \$v3444\ := \$v3443\(0 to 3);
                \$v3438\ := \$v3443\(4 to 35);
                case \$v3444\ is
                when "0010" =>
                  \$1026_i\ := \$v3438\(0 to 31);
                  \$v3442\ := \$arr3237_ptr_take\;
                  if \$v3442\(0) = '1' then
                    \state\ <= q_wait3441;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
                    \state\ <= pause_getI3439;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$369_forever6703194\;
                end case;
              when others =>
                
              end case;
            end if;
          when \$1102_forever6703195\ =>
            \state\ <= \$1102_forever6703195\;
          when \$1114_forever6703224\ =>
            \state\ <= \$1114_forever6703224\;
          when \$1124_forever6703225\ =>
            \state\ <= \$1124_forever6703225\;
          when \$1132_forever6703226\ =>
            \state\ <= \$1132_forever6703226\;
          when \$1137_print_value5913227\ =>
            \$v3481\ := \$1137_print_value5913227_arg\;
            \$v3482\ := \$v3481\(0 to 3);
            \$v3473\ := \$v3481\(4 to 35);
            case \$v3482\ is
            when "0010" =>
              \$1140_t\ := \$v3473\(0 to 31);
              \$v3479\ := "0010" & \$1140_t\;
              \$v3480\ := \$v3479\(0 to 3);
              \$v3474\ := \$v3479\(4 to 35);
              case \$v3480\ is
              when "0010" =>
                \$1026_i\ := \$v3474\(0 to 31);
                \$v3478\ := \$arr3237_ptr_take\;
                if \$v3478\(0) = '1' then
                  \state\ <= q_wait3477;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
                  \state\ <= pause_getI3475;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_rib expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$369_forever6703193\;
              end case;
            when "0000" =>
              \$1137_print_value5913227_result\ := eclat_unit;
              eclat_print_string(of_string("Nil"));
              
              eclat_print_string(of_string("printed tag dfe code\n"));
              
              \$v3471\ := \$1050_loop648_arg\(104 to 139);
              \$v3472\ := \$v3471\(0 to 3);
              \$v3466\ := \$v3471\(4 to 35);
              case \$v3472\ is
              when "0010" =>
                \$1128_t\ := \$v3466\(0 to 31);
                \$v3470\ := \$arr3237_ptr_take\;
                if \$v3470\(0) = '1' then
                  \state\ <= q_wait3469;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1128_t\));
                  \state\ <= pause_getI3467;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_tag_triplet expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1132_forever6703226\;
              end case;
            when "0001" =>
              \$1142_i\ := \$v3473\(0 to 31);
              \$1137_print_value5913227_result\ := eclat_unit;
              eclat_print_int(\$1142_i\);
              
              eclat_print_string(of_string("printed tag dfe code\n"));
              
              \$v3471\ := \$1050_loop648_arg\(104 to 139);
              \$v3472\ := \$v3471\(0 to 3);
              \$v3466\ := \$v3471\(4 to 35);
              case \$v3472\ is
              when "0010" =>
                \$1128_t\ := \$v3466\(0 to 31);
                \$v3470\ := \$arr3237_ptr_take\;
                if \$v3470\(0) = '1' then
                  \state\ <= q_wait3469;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1128_t\));
                  \state\ <= pause_getI3467;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_tag_triplet expected a triplet"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1132_forever6703226\;
              end case;
            when others =>
              
            end case;
          when \$1147_forever6703228\ =>
            \state\ <= \$1147_forever6703228\;
          when \$1164_forever6703229\ =>
            \state\ <= \$1164_forever6703229\;
          when \$1172_forever6703230\ =>
            \state\ <= \$1172_forever6703230\;
          when \$1178_loop6503231\ =>
            \$v3575\ := \$1178_loop6503231_arg\;
            \$v3576\ := \$v3575\(0 to 3);
            \$v3570\ := \$v3575\(4 to 35);
            case \$v3576\ is
            when "0010" =>
              \$1191_t\ := \$v3570\(0 to 31);
              \$v3574\ := \$arr3237_ptr_take\;
              if \$v3574\(0) = '1' then
                \state\ <= q_wait3573;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1191_t\));
                \state\ <= pause_getI3571;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1195_forever6703218\;
            end case;
          when \$1187_forever6703214\ =>
            \state\ <= \$1187_forever6703214\;
          when \$1195_forever6703218\ =>
            \state\ <= \$1195_forever6703218\;
          when \$1229_forever6703232\ =>
            \state\ <= \$1229_forever6703232\;
          when \$1239_forever6703233\ =>
            \state\ <= \$1239_forever6703233\;
          when \$1248_forever6703234\ =>
            \state\ <= \$1248_forever6703234\;
          when \$1260_forever6703235\ =>
            \state\ <= \$1260_forever6703235\;
          when \$1313_forever6703219\ =>
            \state\ <= \$1313_forever6703219\;
          when \$1323_forever6703220\ =>
            \state\ <= \$1323_forever6703220\;
          when \$1332_forever6703221\ =>
            \state\ <= \$1332_forever6703221\;
          when \$1344_forever6703222\ =>
            \state\ <= \$1344_forever6703222\;
          when \$1383_forever6703196\ =>
            \state\ <= \$1383_forever6703196\;
          when \$1398_forever6703197\ =>
            \state\ <= \$1398_forever6703197\;
          when \$369_forever6703193\ =>
            \state\ <= \$369_forever6703193\;
          when \$369_forever6703194\ =>
            \state\ <= \$369_forever6703194\;
          when \$369_forever6703195\ =>
            \state\ <= \$369_forever6703195\;
          when \$369_forever6703216\ =>
            \state\ <= \$369_forever6703216\;
          when \$409_show_rib6123215\ =>
            \$v3542\ := eclat_gt(\$409_show_rib6123215_arg\(68 to 99) & \$409_show_rib6123215_arg\(36 to 67));
            if \$v3542\(0) = '1' then
              \$v3530\ := \$409_show_rib6123215_arg\(0 to 35);
              \$v3531\ := \$v3530\(0 to 3);
              \$v3529\ := \$v3530\(4 to 35);
              case \$v3531\ is
              when "0010" =>
                \$881\ := eclat_true;
                \$v3528\ := \$881\;
                if \$v3528\(0) = '1' then
                  \$409_show_rib6123215_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                  \$1152_k\ := \$1178_loop6503231_result\;
                  \$v3523\ := \$arr3237_ptr_take\;
                  if \$v3523\(0) = '1' then
                    \state\ <= q_wait3522;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                    \state\ <= pause_getI3520;
                  end if;
                else
                  \$v3526\ := \$409_show_rib6123215_arg\(0 to 35);
                  \$v3527\ := \$v3526\(0 to 3);
                  \$v3525\ := \$v3526\(4 to 35);
                  case \$v3527\ is
                  when "0001" =>
                    \$1030_i\ := \$v3525\(0 to 31);
                    \$882\ := \$1030_i\;
                    \$409_show_rib6123215_result\ := eclat_unit;
                    eclat_print_int(\$882\);
                    
                    \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                    \$1152_k\ := \$1178_loop6503231_result\;
                    \$v3523\ := \$arr3237_ptr_take\;
                    if \$v3523\(0) = '1' then
                      \state\ <= q_wait3522;
                    else
                      \$arr3237_ptr_take\(0) := '1';
                      \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                      \state\ <= pause_getI3520;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703195\;
                  end case;
                end if;
              when others =>
                \$881\ := eclat_false;
                \$v3528\ := \$881\;
                if \$v3528\(0) = '1' then
                  \$409_show_rib6123215_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                  \$1152_k\ := \$1178_loop6503231_result\;
                  \$v3523\ := \$arr3237_ptr_take\;
                  if \$v3523\(0) = '1' then
                    \state\ <= q_wait3522;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                    \state\ <= pause_getI3520;
                  end if;
                else
                  \$v3526\ := \$409_show_rib6123215_arg\(0 to 35);
                  \$v3527\ := \$v3526\(0 to 3);
                  \$v3525\ := \$v3526\(4 to 35);
                  case \$v3527\ is
                  when "0001" =>
                    \$1030_i\ := \$v3525\(0 to 31);
                    \$882\ := \$1030_i\;
                    \$409_show_rib6123215_result\ := eclat_unit;
                    eclat_print_int(\$882\);
                    
                    \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                    \$1152_k\ := \$1178_loop6503231_result\;
                    \$v3523\ := \$arr3237_ptr_take\;
                    if \$v3523\(0) = '1' then
                      \state\ <= q_wait3522;
                    else
                      \$arr3237_ptr_take\(0) := '1';
                      \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                      \state\ <= pause_getI3520;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703195\;
                  end case;
                end if;
              end case;
            else
              \$v3540\ := \$409_show_rib6123215_arg\(0 to 35);
              \$v3541\ := \$v3540\(0 to 3);
              \$v3532\ := \$v3540\(4 to 35);
              case \$v3541\ is
              when "0000" =>
                \$409_show_rib6123215_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                \$1152_k\ := \$1178_loop6503231_result\;
                \$v3523\ := \$arr3237_ptr_take\;
                if \$v3523\(0) = '1' then
                  \state\ <= q_wait3522;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                  \state\ <= pause_getI3520;
                end if;
              when "0001" =>
                \$879_i\ := \$v3532\(0 to 31);
                \$409_show_rib6123215_result\ := eclat_unit;
                eclat_print_int(\$879_i\);
                
                \$1178_loop6503231_result\ := \$1178_loop6503231_arg\;
                \$1152_k\ := \$1178_loop6503231_result\;
                \$v3523\ := \$arr3237_ptr_take\;
                if \$v3523\(0) = '1' then
                  \state\ <= q_wait3522;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
                  \state\ <= pause_getI3520;
                end if;
              when "0010" =>
                \$v3538\ := \$409_show_rib6123215_arg\(0 to 35);
                \$v3539\ := \$v3538\(0 to 3);
                \$v3533\ := \$v3538\(4 to 35);
                case \$v3539\ is
                when "0010" =>
                  \$1026_i\ := \$v3533\(0 to 31);
                  \$v3537\ := \$arr3237_ptr_take\;
                  if \$v3537\(0) = '1' then
                    \state\ <= q_wait3536;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
                    \state\ <= pause_getI3534;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$369_forever6703194\;
                end case;
              when others =>
                
              end case;
            end if;
          when \$409_show_rib6123217\ =>
            \$v3567\ := eclat_gt(\$409_show_rib6123217_arg\(68 to 99) & \$409_show_rib6123217_arg\(36 to 67));
            if \$v3567\(0) = '1' then
              \$v3555\ := \$409_show_rib6123217_arg\(0 to 35);
              \$v3556\ := \$v3555\(0 to 3);
              \$v3554\ := \$v3555\(4 to 35);
              case \$v3556\ is
              when "0010" =>
                \$881\ := eclat_true;
                \$v3553\ := \$881\;
                if \$v3553\(0) = '1' then
                  \$409_show_rib6123217_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$v3548\ := \$1178_loop6503231_arg\;
                  \$v3549\ := \$v3548\(0 to 3);
                  \$v3543\ := \$v3548\(4 to 35);
                  case \$v3549\ is
                  when "0010" =>
                    \$977_t\ := \$v3543\(0 to 31);
                    \$v3547\ := \$arr3237_ptr_take\;
                    if \$v3547\(0) = '1' then
                      \state\ <= q_wait3546;
                    else
                      \$arr3237_ptr_take\(0) := '1';
                      \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                      \state\ <= pause_getI3544;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703216\;
                  end case;
                else
                  \$v3551\ := \$409_show_rib6123217_arg\(0 to 35);
                  \$v3552\ := \$v3551\(0 to 3);
                  \$v3550\ := \$v3551\(4 to 35);
                  case \$v3552\ is
                  when "0001" =>
                    \$1030_i\ := \$v3550\(0 to 31);
                    \$882\ := \$1030_i\;
                    \$409_show_rib6123217_result\ := eclat_unit;
                    eclat_print_int(\$882\);
                    
                    \$v3548\ := \$1178_loop6503231_arg\;
                    \$v3549\ := \$v3548\(0 to 3);
                    \$v3543\ := \$v3548\(4 to 35);
                    case \$v3549\ is
                    when "0010" =>
                      \$977_t\ := \$v3543\(0 to 31);
                      \$v3547\ := \$arr3237_ptr_take\;
                      if \$v3547\(0) = '1' then
                        \state\ <= q_wait3546;
                      else
                        \$arr3237_ptr_take\(0) := '1';
                        \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                        \state\ <= pause_getI3544;
                      end if;
                    when others =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \state\ <= \$369_forever6703216\;
                    end case;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703195\;
                  end case;
                end if;
              when others =>
                \$881\ := eclat_false;
                \$v3553\ := \$881\;
                if \$v3553\(0) = '1' then
                  \$409_show_rib6123217_result\ := eclat_unit;
                  eclat_print_string(of_string("[Array]"));
                  
                  \$v3548\ := \$1178_loop6503231_arg\;
                  \$v3549\ := \$v3548\(0 to 3);
                  \$v3543\ := \$v3548\(4 to 35);
                  case \$v3549\ is
                  when "0010" =>
                    \$977_t\ := \$v3543\(0 to 31);
                    \$v3547\ := \$arr3237_ptr_take\;
                    if \$v3547\(0) = '1' then
                      \state\ <= q_wait3546;
                    else
                      \$arr3237_ptr_take\(0) := '1';
                      \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                      \state\ <= pause_getI3544;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703216\;
                  end case;
                else
                  \$v3551\ := \$409_show_rib6123217_arg\(0 to 35);
                  \$v3552\ := \$v3551\(0 to 3);
                  \$v3550\ := \$v3551\(4 to 35);
                  case \$v3552\ is
                  when "0001" =>
                    \$1030_i\ := \$v3550\(0 to 31);
                    \$882\ := \$1030_i\;
                    \$409_show_rib6123217_result\ := eclat_unit;
                    eclat_print_int(\$882\);
                    
                    \$v3548\ := \$1178_loop6503231_arg\;
                    \$v3549\ := \$v3548\(0 to 3);
                    \$v3543\ := \$v3548\(4 to 35);
                    case \$v3549\ is
                    when "0010" =>
                      \$977_t\ := \$v3543\(0 to 31);
                      \$v3547\ := \$arr3237_ptr_take\;
                      if \$v3547\(0) = '1' then
                        \state\ <= q_wait3546;
                      else
                        \$arr3237_ptr_take\(0) := '1';
                        \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                        \state\ <= pause_getI3544;
                      end if;
                    when others =>
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \state\ <= \$369_forever6703216\;
                    end case;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("expected an Integer"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \state\ <= \$369_forever6703195\;
                  end case;
                end if;
              end case;
            else
              \$v3565\ := \$409_show_rib6123217_arg\(0 to 35);
              \$v3566\ := \$v3565\(0 to 3);
              \$v3557\ := \$v3565\(4 to 35);
              case \$v3566\ is
              when "0000" =>
                \$409_show_rib6123217_result\ := eclat_unit;
                eclat_print_string(of_string("Nil"));
                
                \$v3548\ := \$1178_loop6503231_arg\;
                \$v3549\ := \$v3548\(0 to 3);
                \$v3543\ := \$v3548\(4 to 35);
                case \$v3549\ is
                when "0010" =>
                  \$977_t\ := \$v3543\(0 to 31);
                  \$v3547\ := \$arr3237_ptr_take\;
                  if \$v3547\(0) = '1' then
                    \state\ <= q_wait3546;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                    \state\ <= pause_getI3544;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$369_forever6703216\;
                end case;
              when "0001" =>
                \$879_i\ := \$v3557\(0 to 31);
                \$409_show_rib6123217_result\ := eclat_unit;
                eclat_print_int(\$879_i\);
                
                \$v3548\ := \$1178_loop6503231_arg\;
                \$v3549\ := \$v3548\(0 to 3);
                \$v3543\ := \$v3548\(4 to 35);
                case \$v3549\ is
                when "0010" =>
                  \$977_t\ := \$v3543\(0 to 31);
                  \$v3547\ := \$arr3237_ptr_take\;
                  if \$v3547\(0) = '1' then
                    \state\ <= q_wait3546;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
                    \state\ <= pause_getI3544;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$369_forever6703216\;
                end case;
              when "0010" =>
                \$v3563\ := \$409_show_rib6123217_arg\(0 to 35);
                \$v3564\ := \$v3563\(0 to 3);
                \$v3558\ := \$v3563\(4 to 35);
                case \$v3564\ is
                when "0010" =>
                  \$1026_i\ := \$v3558\(0 to 31);
                  \$v3562\ := \$arr3237_ptr_take\;
                  if \$v3562\(0) = '1' then
                    \state\ <= q_wait3561;
                  else
                    \$arr3237_ptr_take\(0) := '1';
                    \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
                    \state\ <= pause_getI3559;
                  end if;
                when others =>
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("get_rib expected a triplet"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \state\ <= \$369_forever6703194\;
                end case;
              when others =>
                
              end case;
            end if;
          when pause_getI3251 =>
            \state\ <= pause_getII3252;
          when pause_getI3259 =>
            \state\ <= pause_getII3260;
          when pause_getI3269 =>
            \state\ <= pause_getII3270;
          when pause_getI3273 =>
            \state\ <= pause_getII3274;
          when pause_getI3277 =>
            \state\ <= pause_getII3278;
          when pause_getI3281 =>
            \state\ <= pause_getII3282;
          when pause_getI3294 =>
            \state\ <= pause_getII3295;
          when pause_getI3306 =>
            \state\ <= pause_getII3307;
          when pause_getI3312 =>
            \state\ <= pause_getII3313;
          when pause_getI3321 =>
            \state\ <= pause_getII3322;
          when pause_getI3327 =>
            \state\ <= pause_getII3328;
          when pause_getI3331 =>
            \state\ <= pause_getII3332;
          when pause_getI3335 =>
            \state\ <= pause_getII3336;
          when pause_getI3350 =>
            \state\ <= pause_getII3351;
          when pause_getI3362 =>
            \state\ <= pause_getII3363;
          when pause_getI3367 =>
            \state\ <= pause_getII3368;
          when pause_getI3372 =>
            \state\ <= pause_getII3373;
          when pause_getI3385 =>
            \state\ <= pause_getII3386;
          when pause_getI3397 =>
            \state\ <= pause_getII3398;
          when pause_getI3403 =>
            \state\ <= pause_getII3404;
          when pause_getI3412 =>
            \state\ <= pause_getII3413;
          when pause_getI3418 =>
            \state\ <= pause_getII3419;
          when pause_getI3422 =>
            \state\ <= pause_getII3423;
          when pause_getI3426 =>
            \state\ <= pause_getII3427;
          when pause_getI3439 =>
            \state\ <= pause_getII3440;
          when pause_getI3448 =>
            \state\ <= pause_getII3449;
          when pause_getI3467 =>
            \state\ <= pause_getII3468;
          when pause_getI3475 =>
            \state\ <= pause_getII3476;
          when pause_getI3484 =>
            \state\ <= pause_getII3485;
          when pause_getI3494 =>
            \state\ <= pause_getII3495;
          when pause_getI3498 =>
            \state\ <= pause_getII3499;
          when pause_getI3507 =>
            \state\ <= pause_getII3508;
          when pause_getI3514 =>
            \state\ <= pause_getII3515;
          when pause_getI3520 =>
            \state\ <= pause_getII3521;
          when pause_getI3534 =>
            \state\ <= pause_getII3535;
          when pause_getI3544 =>
            \state\ <= pause_getII3545;
          when pause_getI3559 =>
            \state\ <= pause_getII3560;
          when pause_getI3571 =>
            \state\ <= pause_getII3572;
          when pause_getI3577 =>
            \state\ <= pause_getII3578;
          when pause_getII3252 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1387\ := \$arr3237_value\;
            \$v3249\ := \$1387\(36 to 71);
            \$v3250\ := \$v3249\(0 to 3);
            \$v3248\ := \$v3249\(4 to 35);
            case \$v3250\ is
            when "0010" =>
              \$1394_i\ := \$v3248\(0 to 31);
              \$1392\ := \$1394_i\;
              \$1391\ := \$1392\ & eclat_sub(\$1046_list_tail618_arg\(32 to 63) & "00000000000000000000000000000001");
              \$1046_list_tail618_arg\ := \$1391\;
              \state\ <= \$1046_list_tail618\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1398_forever6703197\;
            end case;
          when pause_getII3260 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1404\ := \$arr3237_value\;
            \$1402\ := \$1404\(36 to 71);
            \$v3257\ := \$1402\;
            \$v3258\ := \$v3257\(0 to 3);
            \$v3256\ := \$v3257\(4 to 35);
            case \$v3258\ is
            when "0010" =>
              \$1379\ := eclat_true;
              \$v3255\ := \$1379\;
              if \$v3255\(0) = '1' then
                \$v3254\ := \$arr3237_ptr_take\;
                if \$v3254\(0) = '1' then
                  \state\ <= q_wait3253;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1046_list_tail618_arg\(0 to 31)));
                  \state\ <= pause_getI3251;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("list_tail"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1383_forever6703196\;
              end if;
            when others =>
              \$1379\ := eclat_false;
              \$v3255\ := \$1379\;
              if \$v3255\(0) = '1' then
                \$v3254\ := \$arr3237_ptr_take\;
                if \$v3254\(0) = '1' then
                  \state\ <= q_wait3253;
                else
                  \$arr3237_ptr_take\(0) := '1';
                  \$arr3237_ptr\ <= to_integer(unsigned(\$1046_list_tail618_arg\(0 to 31)));
                  \state\ <= pause_getI3251;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("list_tail"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1383_forever6703196\;
              end if;
            end case;
          when pause_getII3270 =>
            \$arr3241_ptr_take\(0) := '0';
            \$1371\ := \$arr3241_value\;
            \$1370\ := \$1371\ & "00000000000000000000000000000001";
            \$1369\ := eclat_add(\$1370\);
            \$v3268\ := \$arr3241_ptr_take\;
            if \$v3268\(0) = '1' then
              \state\ <= q_wait3267;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr_write\ <= 0;
              \$arr3241_write_request\ <= '1';
              \$arr3241_write\ <= \$1369\;
              \state\ <= pause_setI3265;
            end if;
          when pause_getII3274 =>
            \$arr3236_ptr_take\(0) := '0';
            \$1367_c\ := \$arr3236_value\;
            \$v3272\ := \$arr3241_ptr_take\;
            if \$v3272\(0) = '1' then
              \state\ <= q_wait3271;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr\ <= 0;
              \state\ <= pause_getI3269;
            end if;
          when pause_getII3278 =>
            \$arr3241_ptr_take\(0) := '0';
            \$1372\ := \$arr3241_value\;
            \$v3276\ := \$arr3236_ptr_take\;
            if \$v3276\(0) = '1' then
              \state\ <= q_wait3275;
            else
              \$arr3236_ptr_take\(0) := '1';
              \$arr3236_ptr\ <= to_integer(unsigned(\$1372\));
              \state\ <= pause_getI3273;
            end if;
          when pause_getII3282 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1301\ := \$arr3242_value\;
            \$1299\ := "0010" & \$1301\;
            \$1298\ := \$1299\ & eclat_sub(\$1049_rest_loop649_arg\(36 to 67) & "00000000000000000000000000000001");
            \$1049_rest_loop649_arg\ := \$1298\ & \$1049_rest_loop649_arg\(68 to 99) & \$1049_rest_loop649_arg\(100 to 131);
            \state\ <= \$1049_rest_loop649\;
          when pause_getII3295 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1302_i\ := \$arr3242_value\;
            \$v3293\ := \$arr3237_ptr_take\;
            if \$v3293\(0) = '1' then
              \state\ <= q_wait3292;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3289\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1302_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1292\(0 to 35) & \$1049_rest_loop649_arg\(0 to 35) & "0001" & \$v3289\;
              \state\ <= pause_setI3290;
            end if;
          when pause_getII3307 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2830\ := \$arr3237_value\;
            \$1318\ := \$v2830\(36 to 71);
            \$v3303\ := \$1318\;
            \$v3304\ := \$v3303\(0 to 3);
            \$v3302\ := \$v3303\(4 to 35);
            case \$v3304\ is
            when "0010" =>
              \$1319_i\ := \$v3302\(0 to 31);
              \$1317\ := \$1319_i\;
              \$v3301\ := \$arr3238_ptr_take\;
              if \$v3301\(0) = '1' then
                \state\ <= q_wait3300;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr_write\ <= 0;
                \$arr3238_write_request\ <= '1';
                \$arr3238_write\ <= \$1317\;
                \state\ <= pause_setI3298;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1323_forever6703220\;
            end case;
          when pause_getII3313 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1336\ := \$arr3238_value\;
            \$1327\ := "0010" & \$1336\;
            \$v3310\ := \$1327\;
            \$v3311\ := \$v3310\(0 to 3);
            \$v3305\ := \$v3310\(4 to 35);
            case \$v3311\ is
            when "0010" =>
              \$1328_t\ := \$v3305\(0 to 31);
              \$v3309\ := \$arr3237_ptr_take\;
              if \$v3309\(0) = '1' then
                \state\ <= q_wait3308;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1328_t\));
                \state\ <= pause_getI3306;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1332_forever6703221\;
            end case;
          when pause_getII3322 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2834\ := \$arr3237_value\;
            \$1337\ := \$v2834\(36 to 71);
            \$v3318\ := \$1337\;
            \$v3319\ := \$v3318\(0 to 3);
            \$v3317\ := \$v3318\(4 to 35);
            case \$v3319\ is
            when "0010" =>
              \$1309\ := eclat_true;
              \$v3316\ := \$1309\;
              if \$v3316\(0) = '1' then
                \$v3315\ := \$arr3238_ptr_take\;
                if \$v3315\(0) = '1' then
                  \state\ <= q_wait3314;
                else
                  \$arr3238_ptr_take\(0) := '1';
                  \$arr3238_ptr\ <= 0;
                  \state\ <= pause_getI3312;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1313_forever6703219\;
              end if;
            when others =>
              \$1309\ := eclat_false;
              \$v3316\ := \$1309\;
              if \$v3316\(0) = '1' then
                \$v3315\ := \$arr3238_ptr_take\;
                if \$v3315\(0) = '1' then
                  \state\ <= q_wait3314;
                else
                  \$arr3238_ptr_take\(0) := '1';
                  \$arr3238_ptr\ <= 0;
                  \state\ <= pause_getI3312;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1313_forever6703219\;
              end if;
            end case;
          when pause_getII3328 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1348\ := \$arr3238_value\;
            \$1339\ := "0010" & \$1348\;
            \$v3325\ := \$1339\;
            \$v3326\ := \$v3325\(0 to 3);
            \$v3320\ := \$v3325\(4 to 35);
            case \$v3326\ is
            when "0010" =>
              \$1340_t\ := \$v3320\(0 to 31);
              \$v3324\ := \$arr3237_ptr_take\;
              if \$v3324\(0) = '1' then
                \state\ <= q_wait3323;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1340_t\));
                \state\ <= pause_getI3321;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1344_forever6703222\;
            end case;
          when pause_getII3332 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1292\ := \$arr3237_value\;
            \$v3330\ := \$arr3238_ptr_take\;
            if \$v3330\(0) = '1' then
              \state\ <= q_wait3329;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3327;
            end if;
          when pause_getII3336 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1349\ := \$arr3238_value\;
            \$v3334\ := \$arr3237_ptr_take\;
            if \$v3334\(0) = '1' then
              \state\ <= q_wait3333;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1349\));
              \state\ <= pause_getI3331;
            end if;
          when pause_getII3351 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1283\ := \$arr3242_value\;
            \$v3349\ := \$arr3238_ptr_take\;
            if \$v3349\(0) = '1' then
              \state\ <= q_wait3348;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= \$1283\;
              \state\ <= pause_setI3346;
            end if;
          when pause_getII3363 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1285_i\ := \$arr3242_value\;
            \$v3361\ := \$arr3237_ptr_take\;
            if \$v3361\(0) = '1' then
              \state\ <= q_wait3360;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1285_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1284\;
              \state\ <= pause_setI3358;
            end if;
          when pause_getII3368 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1291\ := \$arr3238_value\;
            \$1289\ := "0010" & \$1291\;
            \$v3366\ := "00000000000000000000000000000000";
            \$1284\ := \$1049_rest_loop649_arg\(0 to 35) & \$1289\ & "0001" & \$v3366\;
            \$v3365\ := \$arr3242_ptr_take\;
            if \$v3365\(0) = '1' then
              \state\ <= q_wait3364;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3362;
            end if;
          when pause_getII3373 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1217\ := \$arr3242_value\;
            \$1215\ := "0010" & \$1217\;
            \$1214\ := eclat_sub(\$1050_loop648_arg\(0 to 31) & "00000000000000000000000000000001") & \$1215\;
            \$1050_loop648_arg\ := \$1214\ & \$1050_loop648_arg\(68 to 103) & \$1050_loop648_arg\(104 to 139) & \$1050_loop648_arg\(140 to 171);
            \state\ <= \$1050_loop648\;
          when pause_getII3386 =>
            \$arr3242_ptr_take\(0) := '0';
            \$1218_i\ := \$arr3242_value\;
            \$v3384\ := \$arr3237_ptr_take\;
            if \$v3384\(0) = '1' then
              \state\ <= q_wait3383;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3380\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1218_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1208\(0 to 35) & \$1050_loop648_arg\(32 to 67) & "0001" & \$v3380\;
              \state\ <= pause_setI3381;
            end if;
          when pause_getII3398 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2804\ := \$arr3237_value\;
            \$1234\ := \$v2804\(36 to 71);
            \$v3394\ := \$1234\;
            \$v3395\ := \$v3394\(0 to 3);
            \$v3393\ := \$v3394\(4 to 35);
            case \$v3395\ is
            when "0010" =>
              \$1235_i\ := \$v3393\(0 to 31);
              \$1233\ := \$1235_i\;
              \$v3392\ := \$arr3238_ptr_take\;
              if \$v3392\(0) = '1' then
                \state\ <= q_wait3391;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr_write\ <= 0;
                \$arr3238_write_request\ <= '1';
                \$arr3238_write\ <= \$1233\;
                \state\ <= pause_setI3389;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1239_forever6703233\;
            end case;
          when pause_getII3404 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1252\ := \$arr3238_value\;
            \$1243\ := "0010" & \$1252\;
            \$v3401\ := \$1243\;
            \$v3402\ := \$v3401\(0 to 3);
            \$v3396\ := \$v3401\(4 to 35);
            case \$v3402\ is
            when "0010" =>
              \$1244_t\ := \$v3396\(0 to 31);
              \$v3400\ := \$arr3237_ptr_take\;
              if \$v3400\(0) = '1' then
                \state\ <= q_wait3399;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1244_t\));
                \state\ <= pause_getI3397;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1248_forever6703234\;
            end case;
          when pause_getII3413 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2808\ := \$arr3237_value\;
            \$1253\ := \$v2808\(36 to 71);
            \$v3409\ := \$1253\;
            \$v3410\ := \$v3409\(0 to 3);
            \$v3408\ := \$v3409\(4 to 35);
            case \$v3410\ is
            when "0010" =>
              \$1225\ := eclat_true;
              \$v3407\ := \$1225\;
              if \$v3407\(0) = '1' then
                \$v3406\ := \$arr3238_ptr_take\;
                if \$v3406\(0) = '1' then
                  \state\ <= q_wait3405;
                else
                  \$arr3238_ptr_take\(0) := '1';
                  \$arr3238_ptr\ <= 0;
                  \state\ <= pause_getI3403;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1229_forever6703232\;
              end if;
            when others =>
              \$1225\ := eclat_false;
              \$v3407\ := \$1225\;
              if \$v3407\(0) = '1' then
                \$v3406\ := \$arr3238_ptr_take\;
                if \$v3406\(0) = '1' then
                  \state\ <= q_wait3405;
                else
                  \$arr3238_ptr_take\(0) := '1';
                  \$arr3238_ptr\ <= 0;
                  \state\ <= pause_getI3403;
                end if;
              else
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("get_next_stack"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$1229_forever6703232\;
              end if;
            end case;
          when pause_getII3419 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1264\ := \$arr3238_value\;
            \$1255\ := "0010" & \$1264\;
            \$v3416\ := \$1255\;
            \$v3417\ := \$v3416\(0 to 3);
            \$v3411\ := \$v3416\(4 to 35);
            case \$v3417\ is
            when "0010" =>
              \$1256_t\ := \$v3411\(0 to 31);
              \$v3415\ := \$arr3237_ptr_take\;
              if \$v3415\(0) = '1' then
                \state\ <= q_wait3414;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1256_t\));
                \state\ <= pause_getI3412;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cdr_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1260_forever6703235\;
            end case;
          when pause_getII3423 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1208\ := \$arr3237_value\;
            \$v3421\ := \$arr3238_ptr_take\;
            if \$v3421\(0) = '1' then
              \state\ <= q_wait3420;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3418;
            end if;
          when pause_getII3427 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1265\ := \$arr3238_value\;
            \$v3425\ := \$arr3237_ptr_take\;
            if \$v3425\(0) = '1' then
              \state\ <= q_wait3424;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1265\));
              \state\ <= pause_getI3422;
            end if;
          when pause_getII3440 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3160\ := \$arr3237_value\;
            eclat_print_string(of_string("[ "));
            
            \$1085_show_rib6123223_arg\ := \$v3160\(0 to 35) & \$1085_show_rib6123223_arg\(36 to 67) & eclat_add(\$1085_show_rib6123223_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$1085_show_rib6123223\;
          when pause_getII3449 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1108\ := \$arr3238_value\;
            \$1107\ := "0010" & \$1108\;
            \$1084\ := \$1107\ & "00000000000000000000000000000011" & "00000000000000000000000000000000";
            \$1085_show_rib6123223_arg\ := \$1084\;
            \state\ <= \$1085_show_rib6123223\;
          when pause_getII3468 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2774\ := \$arr3237_value\;
            \$1119\ := \$v2774\(72 to 107);
            \$v3464\ := \$1119\;
            \$v3465\ := \$v3464\(0 to 3);
            \$v3463\ := \$v3464\(4 to 35);
            case \$v3465\ is
            when "0010" =>
              \$1120_i\ := \$v3463\(0 to 31);
              \$1118\ := \$1120_i\;
              \$v3462\ := \$arr3239_ptr_take\;
              if \$v3462\(0) = '1' then
                \state\ <= q_wait3461;
              else
                \$arr3239_ptr_take\(0) := '1';
                \$arr3239_ptr_write\ <= 0;
                \$arr3239_write_request\ <= '1';
                \$arr3239_write\ <= \$1118\;
                \state\ <= pause_setI3459;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1124_forever6703225\;
            end case;
          when pause_getII3476 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3173\ := \$arr3237_value\;
            eclat_print_string(of_string("["));
            
            \$1137_print_value5913227_arg\ := \$v3173\(0 to 35);
            \state\ <= \$1137_print_value5913227\;
          when pause_getII3485 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2778\ := \$arr3237_value\;
            \$1136\ := \$v2778\(72 to 107);
            \$1137_print_value5913227_arg\ := \$1136\;
            \state\ <= \$1137_print_value5913227\;
          when pause_getII3495 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1206\ := \$arr3238_value\;
            \$1205\ := "0010" & \$1206\;
            \$1204\ := \$1205\ & \$1200\(36 to 71) & \$1050_loop648_arg\(68 to 103);
            \$v3493\ := \$arr3237_ptr_take\;
            if \$v3493\(0) = '1' then
              \state\ <= q_wait3492;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1204\;
              \state\ <= pause_setI3490;
            end if;
          when pause_getII3499 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1200\ := \$arr3237_value\;
            \$v3497\ := \$arr3238_ptr_take\;
            if \$v3497\(0) = '1' then
              \state\ <= q_wait3496;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3494;
            end if;
          when pause_getII3508 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2783\ := \$arr3237_value\;
            \$1159\ := \$v2783\(72 to 107);
            \$1157\ := \$1158\ & \$1153\(36 to 71) & \$1159\;
            \$v3505\ := \$arr3237_ptr_take\;
            if \$v3505\(0) = '1' then
              \state\ <= q_wait3504;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1157\;
              \state\ <= pause_setI3502;
            end if;
          when pause_getII3515 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2787\ := \$arr3237_value\;
            \$1158\ := \$v2787\(0 to 35);
            \$v3511\ := \$1152_k\;
            \$v3512\ := \$v3511\(0 to 3);
            \$v3506\ := \$v3511\(4 to 35);
            case \$v3512\ is
            when "0010" =>
              \$1160_t\ := \$v3506\(0 to 31);
              \$v3510\ := \$arr3237_ptr_take\;
              if \$v3510\(0) = '1' then
                \state\ <= q_wait3509;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1160_t\));
                \state\ <= pause_getI3507;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1164_forever6703229\;
            end case;
          when pause_getII3521 =>
            \$arr3237_ptr_take\(0) := '0';
            \$1153\ := \$arr3237_value\;
            \$v3518\ := \$1152_k\;
            \$v3519\ := \$v3518\(0 to 3);
            \$v3513\ := \$v3518\(4 to 35);
            case \$v3519\ is
            when "0010" =>
              \$1168_t\ := \$v3513\(0 to 31);
              \$v3517\ := \$arr3237_ptr_take\;
              if \$v3517\(0) = '1' then
                \state\ <= q_wait3516;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1168_t\));
                \state\ <= pause_getI3514;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_car_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1172_forever6703230\;
            end case;
          when pause_getII3535 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3160\ := \$arr3237_value\;
            eclat_print_string(of_string("[ "));
            
            \$409_show_rib6123215_arg\ := \$v3160\(0 to 35) & \$409_show_rib6123215_arg\(36 to 67) & eclat_add(\$409_show_rib6123215_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$409_show_rib6123215\;
          when pause_getII3545 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2843\ := \$arr3237_value\;
            \$v405\ := \$v2843\(36 to 71);
            \$1178_loop6503231_arg\ := \$v405\;
            \state\ <= \$1178_loop6503231\;
          when pause_getII3560 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3160\ := \$arr3237_value\;
            eclat_print_string(of_string("[ "));
            
            \$409_show_rib6123217_arg\ := \$v3160\(0 to 35) & \$409_show_rib6123217_arg\(36 to 67) & eclat_add(\$409_show_rib6123217_arg\(68 to 99) & "00000000000000000000000000000001");
            \state\ <= \$409_show_rib6123217\;
          when pause_getII3572 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v2847\ := \$arr3237_value\;
            \$1181_tag\ := \$v2847\(72 to 107);
            \$v3568\ := \$1181_tag\;
            \$v3569\ := \$v3568\(0 to 3);
            \$v3524\ := \$v3568\(4 to 35);
            case \$v3569\ is
            when "0010" =>
              \$409_show_rib6123215_arg\ := \$1178_loop6503231_arg\ & "00000000000000000000000000000101" & "00000000000000000000000000000000";
              \state\ <= \$409_show_rib6123215\;
            when "0001" =>
              \$409_show_rib6123217_arg\ := \$1178_loop6503231_arg\ & "00000000000000000000000000000101" & "00000000000000000000000000000000";
              \state\ <= \$409_show_rib6123217\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_cont 2"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1187_forever6703214\;
            end case;
          when pause_getII3578 =>
            \$arr3238_ptr_take\(0) := '0';
            \$1199\ := \$arr3238_value\;
            \$1177\ := "0010" & \$1199\;
            \$1178_loop6503231_arg\ := \$1177\;
            \state\ <= \$1178_loop6503231\;
          when pause_setI3265 =>
            \$arr3241_write_request\ <= '0';
            \state\ <= pause_setII3266;
          when pause_setI3285 =>
            \$arr3242_write_request\ <= '0';
            \state\ <= pause_setII3286;
          when pause_setI3290 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3291;
          when pause_setI3298 =>
            \$arr3238_write_request\ <= '0';
            \state\ <= pause_setII3299;
          when pause_setI3342 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3343;
          when pause_setI3346 =>
            \$arr3238_write_request\ <= '0';
            \state\ <= pause_setII3347;
          when pause_setI3354 =>
            \$arr3242_write_request\ <= '0';
            \state\ <= pause_setII3355;
          when pause_setI3358 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3359;
          when pause_setI3376 =>
            \$arr3242_write_request\ <= '0';
            \state\ <= pause_setII3377;
          when pause_setI3381 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3382;
          when pause_setI3389 =>
            \$arr3238_write_request\ <= '0';
            \state\ <= pause_setII3390;
          when pause_setI3452 =>
            \$arr3238_write_request\ <= '0';
            \state\ <= pause_setII3453;
          when pause_setI3459 =>
            \$arr3239_write_request\ <= '0';
            \state\ <= pause_setII3460;
          when pause_setI3490 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3491;
          when pause_setI3502 =>
            \$arr3237_write_request\ <= '0';
            \state\ <= pause_setII3503;
          when pause_setI3586 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3587;
          when pause_setI3590 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3591;
          when pause_setI3594 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3595;
          when pause_setI3598 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3599;
          when pause_setI3602 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3603;
          when pause_setI3606 =>
            \$arr3243_write_request\ <= '0';
            \state\ <= pause_setII3607;
          when pause_setI3610 =>
            \$arr3242_write_request\ <= '0';
            \state\ <= pause_setII3611;
          when pause_setI3614 =>
            \$arr3241_write_request\ <= '0';
            \state\ <= pause_setII3615;
          when pause_setI3618 =>
            \$arr3240_write_request\ <= '0';
            \state\ <= pause_setII3619;
          when pause_setI3622 =>
            \$arr3238_write_request\ <= '0';
            \state\ <= pause_setII3623;
          when pause_setI3626 =>
            \$arr3239_write_request\ <= '0';
            \state\ <= pause_setII3627;
          when pause_setII3266 =>
            \$arr3241_ptr_take\(0) := '0';
            \$1365\ := \$1367_c\;
            \$1364\ := \$1365\ & X"000000" & X"23";
            \$1362_x\ := eclat_sub(\$1364\);
            \$1352_x\ := eclat_if(eclat_lt(\$1362_x\ & "00000000000000000000000000000000") & X"000000" & X"39" & \$1362_x\);
            \$v3264\ := eclat_lt(\$1352_x\ & X"000000" & X"2e");
            if \$v3264\(0) = '1' then
              \state\ <= \$1047_get_int621\;
            else
              \$1047_get_int621_arg\ := eclat_sub(eclat_add(eclat_mult(\$1047_get_int621_arg\ & X"000000" & X"2e") & \$1352_x\) & X"000000" & X"2e");
              \state\ <= \$1047_get_int621\;
            end if;
          when pause_setII3286 =>
            \$arr3242_ptr_take\(0) := '0';
            \$v3284\ := \$arr3242_ptr_take\;
            if \$v3284\(0) = '1' then
              \state\ <= q_wait3283;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3281;
            end if;
          when pause_setII3291 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3288\ := \$arr3242_ptr_take\;
            if \$v3288\(0) = '1' then
              \state\ <= q_wait3287;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1302_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3285;
            end if;
          when pause_setII3299 =>
            \$arr3238_ptr_take\(0) := '0';
            \$v3297\ := \$arr3242_ptr_take\;
            if \$v3297\(0) = '1' then
              \state\ <= q_wait3296;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3294;
            end if;
          when pause_setII3343 =>
            \$arr3237_ptr_take\(0) := '0';
            \state\ <= \$1049_rest_loop649\;
          when pause_setII3347 =>
            \$arr3238_ptr_take\(0) := '0';
            \$v3345\ := \$arr3237_ptr_take\;
            if \$v3345\(0) = '1' then
              \state\ <= q_wait3344;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3339\ := eclat_add(\$1049_rest_loop649_arg\(100 to 131) & "00000000000000000000000000000001");
              \$v3340\ := "00000000000000000000000000000000";
              \$v3341\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1049_rest_loop649_arg\(68 to 99)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= "0001" & \$v3339\ & "0001" & \$v3340\ & "0001" & \$v3341\;
              \state\ <= pause_setI3342;
            end if;
          when pause_setII3355 =>
            \$arr3242_ptr_take\(0) := '0';
            \$v3353\ := \$arr3242_ptr_take\;
            if \$v3353\(0) = '1' then
              \state\ <= q_wait3352;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3350;
            end if;
          when pause_setII3359 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3357\ := \$arr3242_ptr_take\;
            if \$v3357\(0) = '1' then
              \state\ <= q_wait3356;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1285_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3354;
            end if;
          when pause_setII3377 =>
            \$arr3242_ptr_take\(0) := '0';
            \$v3375\ := \$arr3242_ptr_take\;
            if \$v3375\(0) = '1' then
              \state\ <= q_wait3374;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3372;
            end if;
          when pause_setII3382 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3379\ := \$arr3242_ptr_take\;
            if \$v3379\(0) = '1' then
              \state\ <= q_wait3378;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1218_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3376;
            end if;
          when pause_setII3390 =>
            \$arr3238_ptr_take\(0) := '0';
            \$v3388\ := \$arr3242_ptr_take\;
            if \$v3388\(0) = '1' then
              \state\ <= q_wait3387;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3385;
            end if;
          when pause_setII3453 =>
            \$arr3238_ptr_take\(0) := '0';
            \$v3451\ := \$arr3238_ptr_take\;
            if \$v3451\(0) = '1' then
              \state\ <= q_wait3450;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3448;
            end if;
          when pause_setII3460 =>
            \$arr3239_ptr_take\(0) := '0';
            \$v3457\ := \$1050_loop648_arg\(32 to 67);
            \$v3458\ := \$v3457\(0 to 3);
            \$v3456\ := \$v3457\(4 to 35);
            case \$v3458\ is
            when "0010" =>
              \$1110_i\ := \$v3456\(0 to 31);
              \$1109\ := \$1110_i\;
              \$v3455\ := \$arr3238_ptr_take\;
              if \$v3455\(0) = '1' then
                \state\ <= q_wait3454;
              else
                \$arr3238_ptr_take\(0) := '1';
                \$arr3238_ptr_write\ <= 0;
                \$arr3238_write_request\ <= '1';
                \$arr3238_write\ <= \$1109\;
                \state\ <= pause_setI3452;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("expected a triplet 1"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1114_forever6703224\;
            end case;
          when pause_setII3491 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3488\ := \$1050_loop648_arg\(104 to 139);
            \$v3489\ := \$v3488\(0 to 3);
            \$v3483\ := \$v3488\(4 to 35);
            case \$v3489\ is
            when "0010" =>
              \$1143_t\ := \$v3483\(0 to 31);
              \$v3487\ := \$arr3237_ptr_take\;
              if \$v3487\(0) = '1' then
                \state\ <= q_wait3486;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1143_t\));
                \state\ <= pause_getI3484;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1147_forever6703228\;
            end case;
          when pause_setII3503 =>
            \$arr3237_ptr_take\(0) := '0';
            \$v3488\ := \$1050_loop648_arg\(104 to 139);
            \$v3489\ := \$v3488\(0 to 3);
            \$v3483\ := \$v3488\(4 to 35);
            case \$v3489\ is
            when "0010" =>
              \$1143_t\ := \$v3483\(0 to 31);
              \$v3487\ := \$arr3237_ptr_take\;
              if \$v3487\(0) = '1' then
                \state\ <= q_wait3486;
              else
                \$arr3237_ptr_take\(0) := '1';
                \$arr3237_ptr\ <= to_integer(unsigned(\$1143_t\));
                \state\ <= pause_getI3484;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("get_tag_triplet expected a triplet"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$1147_forever6703228\;
            end case;
          when pause_setII3587 =>
            \$arr3243_ptr_take\(0) := '0';
            eclat_print_string(of_string("Compilation reussi, pas de bug dans la syntaxe "));
            
            result3244 := eclat_unit;
            eclat_print_newline(eclat_unit);
            
            rdy3245 := eclat_true;
            \state\ <= compute3246;
          when pause_setII3591 =>
            \$arr3243_ptr_take\(0) := '0';
            \$v3589\ := \$arr3243_ptr_take\;
            if \$v3589\(0) = '1' then
              \state\ <= q_wait3588;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 5;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI3586;
            end if;
          when pause_setII3595 =>
            \$arr3243_ptr_take\(0) := '0';
            \$v3593\ := \$arr3243_ptr_take\;
            if \$v3593\(0) = '1' then
              \state\ <= q_wait3592;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 4;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI3590;
            end if;
          when pause_setII3599 =>
            \$arr3243_ptr_take\(0) := '0';
            \$v3597\ := \$arr3243_ptr_take\;
            if \$v3597\(0) = '1' then
              \state\ <= q_wait3596;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 3;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI3594;
            end if;
          when pause_setII3603 =>
            \$arr3243_ptr_take\(0) := '0';
            \$v3601\ := \$arr3243_ptr_take\;
            if \$v3601\(0) = '1' then
              \state\ <= q_wait3600;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 2;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI3598;
            end if;
          when pause_setII3607 =>
            \$arr3243_ptr_take\(0) := '0';
            \$v3605\ := \$arr3243_ptr_take\;
            if \$v3605\(0) = '1' then
              \state\ <= q_wait3604;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 1;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI3602;
            end if;
          when pause_setII3611 =>
            \$arr3242_ptr_take\(0) := '0';
            \$v3609\ := \$arr3243_ptr_take\;
            if \$v3609\(0) = '1' then
              \state\ <= q_wait3608;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 0;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= X"000000" & X"14";
              \state\ <= pause_setI3606;
            end if;
          when pause_setII3615 =>
            \$arr3241_ptr_take\(0) := '0';
            \$v3613\ := \$arr3242_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3610;
            end if;
          when pause_setII3619 =>
            \$arr3240_ptr_take\(0) := '0';
            \$v3617\ := \$arr3241_ptr_take\;
            if \$v3617\(0) = '1' then
              \state\ <= q_wait3616;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr_write\ <= 0;
              \$arr3241_write_request\ <= '1';
              \$arr3241_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI3614;
            end if;
          when pause_setII3623 =>
            \$arr3238_ptr_take\(0) := '0';
            \$v3621\ := \$arr3240_ptr_take\;
            if \$v3621\(0) = '1' then
              \state\ <= q_wait3620;
            else
              \$arr3240_ptr_take\(0) := '1';
              \$arr3240_ptr_write\ <= 0;
              \$arr3240_write_request\ <= '1';
              \$arr3240_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3618;
            end if;
          when pause_setII3627 =>
            \$arr3239_ptr_take\(0) := '0';
            \$v3625\ := \$arr3238_ptr_take\;
            if \$v3625\(0) = '1' then
              \state\ <= q_wait3624;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI3622;
            end if;
          when q_wait3253 =>
            \$v3254\ := \$arr3237_ptr_take\;
            if \$v3254\(0) = '1' then
              \state\ <= q_wait3253;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1046_list_tail618_arg\(0 to 31)));
              \state\ <= pause_getI3251;
            end if;
          when q_wait3261 =>
            \$v3262\ := \$arr3237_ptr_take\;
            if \$v3262\(0) = '1' then
              \state\ <= q_wait3261;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1046_list_tail618_arg\(0 to 31)));
              \state\ <= pause_getI3259;
            end if;
          when q_wait3267 =>
            \$v3268\ := \$arr3241_ptr_take\;
            if \$v3268\(0) = '1' then
              \state\ <= q_wait3267;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr_write\ <= 0;
              \$arr3241_write_request\ <= '1';
              \$arr3241_write\ <= \$1369\;
              \state\ <= pause_setI3265;
            end if;
          when q_wait3271 =>
            \$v3272\ := \$arr3241_ptr_take\;
            if \$v3272\(0) = '1' then
              \state\ <= q_wait3271;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr\ <= 0;
              \state\ <= pause_getI3269;
            end if;
          when q_wait3275 =>
            \$v3276\ := \$arr3236_ptr_take\;
            if \$v3276\(0) = '1' then
              \state\ <= q_wait3275;
            else
              \$arr3236_ptr_take\(0) := '1';
              \$arr3236_ptr\ <= to_integer(unsigned(\$1372\));
              \state\ <= pause_getI3273;
            end if;
          when q_wait3279 =>
            \$v3280\ := \$arr3241_ptr_take\;
            if \$v3280\(0) = '1' then
              \state\ <= q_wait3279;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr\ <= 0;
              \state\ <= pause_getI3277;
            end if;
          when q_wait3283 =>
            \$v3284\ := \$arr3242_ptr_take\;
            if \$v3284\(0) = '1' then
              \state\ <= q_wait3283;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3281;
            end if;
          when q_wait3287 =>
            \$v3288\ := \$arr3242_ptr_take\;
            if \$v3288\(0) = '1' then
              \state\ <= q_wait3287;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1302_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3285;
            end if;
          when q_wait3292 =>
            \$v3293\ := \$arr3237_ptr_take\;
            if \$v3293\(0) = '1' then
              \state\ <= q_wait3292;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3289\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1302_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1292\(0 to 35) & \$1049_rest_loop649_arg\(0 to 35) & "0001" & \$v3289\;
              \state\ <= pause_setI3290;
            end if;
          when q_wait3296 =>
            \$v3297\ := \$arr3242_ptr_take\;
            if \$v3297\(0) = '1' then
              \state\ <= q_wait3296;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3294;
            end if;
          when q_wait3300 =>
            \$v3301\ := \$arr3238_ptr_take\;
            if \$v3301\(0) = '1' then
              \state\ <= q_wait3300;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= \$1317\;
              \state\ <= pause_setI3298;
            end if;
          when q_wait3308 =>
            \$v3309\ := \$arr3237_ptr_take\;
            if \$v3309\(0) = '1' then
              \state\ <= q_wait3308;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1328_t\));
              \state\ <= pause_getI3306;
            end if;
          when q_wait3314 =>
            \$v3315\ := \$arr3238_ptr_take\;
            if \$v3315\(0) = '1' then
              \state\ <= q_wait3314;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3312;
            end if;
          when q_wait3323 =>
            \$v3324\ := \$arr3237_ptr_take\;
            if \$v3324\(0) = '1' then
              \state\ <= q_wait3323;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1340_t\));
              \state\ <= pause_getI3321;
            end if;
          when q_wait3329 =>
            \$v3330\ := \$arr3238_ptr_take\;
            if \$v3330\(0) = '1' then
              \state\ <= q_wait3329;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3327;
            end if;
          when q_wait3333 =>
            \$v3334\ := \$arr3237_ptr_take\;
            if \$v3334\(0) = '1' then
              \state\ <= q_wait3333;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1349\));
              \state\ <= pause_getI3331;
            end if;
          when q_wait3337 =>
            \$v3338\ := \$arr3238_ptr_take\;
            if \$v3338\(0) = '1' then
              \state\ <= q_wait3337;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3335;
            end if;
          when q_wait3344 =>
            \$v3345\ := \$arr3237_ptr_take\;
            if \$v3345\(0) = '1' then
              \state\ <= q_wait3344;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3339\ := eclat_add(\$1049_rest_loop649_arg\(100 to 131) & "00000000000000000000000000000001");
              \$v3340\ := "00000000000000000000000000000000";
              \$v3341\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1049_rest_loop649_arg\(68 to 99)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= "0001" & \$v3339\ & "0001" & \$v3340\ & "0001" & \$v3341\;
              \state\ <= pause_setI3342;
            end if;
          when q_wait3348 =>
            \$v3349\ := \$arr3238_ptr_take\;
            if \$v3349\(0) = '1' then
              \state\ <= q_wait3348;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= \$1283\;
              \state\ <= pause_setI3346;
            end if;
          when q_wait3352 =>
            \$v3353\ := \$arr3242_ptr_take\;
            if \$v3353\(0) = '1' then
              \state\ <= q_wait3352;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3350;
            end if;
          when q_wait3356 =>
            \$v3357\ := \$arr3242_ptr_take\;
            if \$v3357\(0) = '1' then
              \state\ <= q_wait3356;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1285_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3354;
            end if;
          when q_wait3360 =>
            \$v3361\ := \$arr3237_ptr_take\;
            if \$v3361\(0) = '1' then
              \state\ <= q_wait3360;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1285_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1284\;
              \state\ <= pause_setI3358;
            end if;
          when q_wait3364 =>
            \$v3365\ := \$arr3242_ptr_take\;
            if \$v3365\(0) = '1' then
              \state\ <= q_wait3364;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3362;
            end if;
          when q_wait3369 =>
            \$v3370\ := \$arr3238_ptr_take\;
            if \$v3370\(0) = '1' then
              \state\ <= q_wait3369;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3367;
            end if;
          when q_wait3374 =>
            \$v3375\ := \$arr3242_ptr_take\;
            if \$v3375\(0) = '1' then
              \state\ <= q_wait3374;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3372;
            end if;
          when q_wait3378 =>
            \$v3379\ := \$arr3242_ptr_take\;
            if \$v3379\(0) = '1' then
              \state\ <= q_wait3378;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub(\$1218_i\ & "00000000000000000000000000000001");
              \state\ <= pause_setI3376;
            end if;
          when q_wait3383 =>
            \$v3384\ := \$arr3237_ptr_take\;
            if \$v3384\(0) = '1' then
              \state\ <= q_wait3383;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$v3380\ := "00000000000000000000000000000000";
              \$arr3237_ptr_write\ <= to_integer(unsigned(eclat_sub(\$1218_i\ & "00000000000000000000000000000001")));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1208\(0 to 35) & \$1050_loop648_arg\(32 to 67) & "0001" & \$v3380\;
              \state\ <= pause_setI3381;
            end if;
          when q_wait3387 =>
            \$v3388\ := \$arr3242_ptr_take\;
            if \$v3388\(0) = '1' then
              \state\ <= q_wait3387;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr\ <= 0;
              \state\ <= pause_getI3385;
            end if;
          when q_wait3391 =>
            \$v3392\ := \$arr3238_ptr_take\;
            if \$v3392\(0) = '1' then
              \state\ <= q_wait3391;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= \$1233\;
              \state\ <= pause_setI3389;
            end if;
          when q_wait3399 =>
            \$v3400\ := \$arr3237_ptr_take\;
            if \$v3400\(0) = '1' then
              \state\ <= q_wait3399;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1244_t\));
              \state\ <= pause_getI3397;
            end if;
          when q_wait3405 =>
            \$v3406\ := \$arr3238_ptr_take\;
            if \$v3406\(0) = '1' then
              \state\ <= q_wait3405;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3403;
            end if;
          when q_wait3414 =>
            \$v3415\ := \$arr3237_ptr_take\;
            if \$v3415\(0) = '1' then
              \state\ <= q_wait3414;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1256_t\));
              \state\ <= pause_getI3412;
            end if;
          when q_wait3420 =>
            \$v3421\ := \$arr3238_ptr_take\;
            if \$v3421\(0) = '1' then
              \state\ <= q_wait3420;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3418;
            end if;
          when q_wait3424 =>
            \$v3425\ := \$arr3237_ptr_take\;
            if \$v3425\(0) = '1' then
              \state\ <= q_wait3424;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1265\));
              \state\ <= pause_getI3422;
            end if;
          when q_wait3428 =>
            \$v3429\ := \$arr3238_ptr_take\;
            if \$v3429\(0) = '1' then
              \state\ <= q_wait3428;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3426;
            end if;
          when q_wait3441 =>
            \$v3442\ := \$arr3237_ptr_take\;
            if \$v3442\(0) = '1' then
              \state\ <= q_wait3441;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
              \state\ <= pause_getI3439;
            end if;
          when q_wait3450 =>
            \$v3451\ := \$arr3238_ptr_take\;
            if \$v3451\(0) = '1' then
              \state\ <= q_wait3450;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3448;
            end if;
          when q_wait3454 =>
            \$v3455\ := \$arr3238_ptr_take\;
            if \$v3455\(0) = '1' then
              \state\ <= q_wait3454;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= \$1109\;
              \state\ <= pause_setI3452;
            end if;
          when q_wait3461 =>
            \$v3462\ := \$arr3239_ptr_take\;
            if \$v3462\(0) = '1' then
              \state\ <= q_wait3461;
            else
              \$arr3239_ptr_take\(0) := '1';
              \$arr3239_ptr_write\ <= 0;
              \$arr3239_write_request\ <= '1';
              \$arr3239_write\ <= \$1118\;
              \state\ <= pause_setI3459;
            end if;
          when q_wait3469 =>
            \$v3470\ := \$arr3237_ptr_take\;
            if \$v3470\(0) = '1' then
              \state\ <= q_wait3469;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1128_t\));
              \state\ <= pause_getI3467;
            end if;
          when q_wait3477 =>
            \$v3478\ := \$arr3237_ptr_take\;
            if \$v3478\(0) = '1' then
              \state\ <= q_wait3477;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
              \state\ <= pause_getI3475;
            end if;
          when q_wait3486 =>
            \$v3487\ := \$arr3237_ptr_take\;
            if \$v3487\(0) = '1' then
              \state\ <= q_wait3486;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1143_t\));
              \state\ <= pause_getI3484;
            end if;
          when q_wait3492 =>
            \$v3493\ := \$arr3237_ptr_take\;
            if \$v3493\(0) = '1' then
              \state\ <= q_wait3492;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1204\;
              \state\ <= pause_setI3490;
            end if;
          when q_wait3496 =>
            \$v3497\ := \$arr3238_ptr_take\;
            if \$v3497\(0) = '1' then
              \state\ <= q_wait3496;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3494;
            end if;
          when q_wait3500 =>
            \$v3501\ := \$arr3237_ptr_take\;
            if \$v3501\(0) = '1' then
              \state\ <= q_wait3500;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \state\ <= pause_getI3498;
            end if;
          when q_wait3504 =>
            \$v3505\ := \$arr3237_ptr_take\;
            if \$v3505\(0) = '1' then
              \state\ <= q_wait3504;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr_write\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \$arr3237_write_request\ <= '1';
              \$arr3237_write\ <= \$1157\;
              \state\ <= pause_setI3502;
            end if;
          when q_wait3509 =>
            \$v3510\ := \$arr3237_ptr_take\;
            if \$v3510\(0) = '1' then
              \state\ <= q_wait3509;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1160_t\));
              \state\ <= pause_getI3507;
            end if;
          when q_wait3516 =>
            \$v3517\ := \$arr3237_ptr_take\;
            if \$v3517\(0) = '1' then
              \state\ <= q_wait3516;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1168_t\));
              \state\ <= pause_getI3514;
            end if;
          when q_wait3522 =>
            \$v3523\ := \$arr3237_ptr_take\;
            if \$v3523\(0) = '1' then
              \state\ <= q_wait3522;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1050_loop648_arg\(140 to 171)));
              \state\ <= pause_getI3520;
            end if;
          when q_wait3536 =>
            \$v3537\ := \$arr3237_ptr_take\;
            if \$v3537\(0) = '1' then
              \state\ <= q_wait3536;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
              \state\ <= pause_getI3534;
            end if;
          when q_wait3546 =>
            \$v3547\ := \$arr3237_ptr_take\;
            if \$v3547\(0) = '1' then
              \state\ <= q_wait3546;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$977_t\));
              \state\ <= pause_getI3544;
            end if;
          when q_wait3561 =>
            \$v3562\ := \$arr3237_ptr_take\;
            if \$v3562\(0) = '1' then
              \state\ <= q_wait3561;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1026_i\));
              \state\ <= pause_getI3559;
            end if;
          when q_wait3573 =>
            \$v3574\ := \$arr3237_ptr_take\;
            if \$v3574\(0) = '1' then
              \state\ <= q_wait3573;
            else
              \$arr3237_ptr_take\(0) := '1';
              \$arr3237_ptr\ <= to_integer(unsigned(\$1191_t\));
              \state\ <= pause_getI3571;
            end if;
          when q_wait3579 =>
            \$v3580\ := \$arr3238_ptr_take\;
            if \$v3580\(0) = '1' then
              \state\ <= q_wait3579;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr\ <= 0;
              \state\ <= pause_getI3577;
            end if;
          when q_wait3588 =>
            \$v3589\ := \$arr3243_ptr_take\;
            if \$v3589\(0) = '1' then
              \state\ <= q_wait3588;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 5;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000000100";
              \state\ <= pause_setI3586;
            end if;
          when q_wait3592 =>
            \$v3593\ := \$arr3243_ptr_take\;
            if \$v3593\(0) = '1' then
              \state\ <= q_wait3592;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 4;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000001011";
              \state\ <= pause_setI3590;
            end if;
          when q_wait3596 =>
            \$v3597\ := \$arr3243_ptr_take\;
            if \$v3597\(0) = '1' then
              \state\ <= q_wait3596;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 3;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000001010";
              \state\ <= pause_setI3594;
            end if;
          when q_wait3600 =>
            \$v3601\ := \$arr3243_ptr_take\;
            if \$v3601\(0) = '1' then
              \state\ <= q_wait3600;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 2;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI3598;
            end if;
          when q_wait3604 =>
            \$v3605\ := \$arr3243_ptr_take\;
            if \$v3605\(0) = '1' then
              \state\ <= q_wait3604;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 1;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= X"000000" & X"1e";
              \state\ <= pause_setI3602;
            end if;
          when q_wait3608 =>
            \$v3609\ := \$arr3243_ptr_take\;
            if \$v3609\(0) = '1' then
              \state\ <= q_wait3608;
            else
              \$arr3243_ptr_take\(0) := '1';
              \$arr3243_ptr_write\ <= 0;
              \$arr3243_write_request\ <= '1';
              \$arr3243_write\ <= X"000000" & X"14";
              \state\ <= pause_setI3606;
            end if;
          when q_wait3612 =>
            \$v3613\ := \$arr3242_ptr_take\;
            if \$v3613\(0) = '1' then
              \state\ <= q_wait3612;
            else
              \$arr3242_ptr_take\(0) := '1';
              \$arr3242_ptr_write\ <= 0;
              \$arr3242_write_request\ <= '1';
              \$arr3242_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3610;
            end if;
          when q_wait3616 =>
            \$v3617\ := \$arr3241_ptr_take\;
            if \$v3617\(0) = '1' then
              \state\ <= q_wait3616;
            else
              \$arr3241_ptr_take\(0) := '1';
              \$arr3241_ptr_write\ <= 0;
              \$arr3241_write_request\ <= '1';
              \$arr3241_write\ <= "00000000000000000000000000000000";
              \state\ <= pause_setI3614;
            end if;
          when q_wait3620 =>
            \$v3621\ := \$arr3240_ptr_take\;
            if \$v3621\(0) = '1' then
              \state\ <= q_wait3620;
            else
              \$arr3240_ptr_take\(0) := '1';
              \$arr3240_ptr_write\ <= 0;
              \$arr3240_write_request\ <= '1';
              \$arr3240_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3618;
            end if;
          when q_wait3624 =>
            \$v3625\ := \$arr3238_ptr_take\;
            if \$v3625\(0) = '1' then
              \state\ <= q_wait3624;
            else
              \$arr3238_ptr_take\(0) := '1';
              \$arr3238_ptr_write\ <= 0;
              \$arr3238_write_request\ <= '1';
              \$arr3238_write\ <= X"0000" & X"2328";
              \state\ <= pause_setI3622;
            end if;
          when q_wait3628 =>
            \$v3629\ := \$arr3239_ptr_take\;
            if \$v3629\(0) = '1' then
              \state\ <= q_wait3628;
            else
              \$arr3239_ptr_take\(0) := '1';
              \$arr3239_ptr_write\ <= 0;
              \$arr3239_write_request\ <= '1';
              \$arr3239_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3626;
            end if;
          when compute3246 =>
            rdy3245 := eclat_false;
            \$v3629\ := \$arr3239_ptr_take\;
            if \$v3629\(0) = '1' then
              \state\ <= q_wait3628;
            else
              \$arr3239_ptr_take\(0) := '1';
              \$arr3239_ptr_write\ <= 0;
              \$arr3239_write_request\ <= '1';
              \$arr3239_write\ <= eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001");
              \state\ <= pause_setI3626;
            end if;
          end case;
          
          result <= result3244;
          rdy <= rdy3245;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
